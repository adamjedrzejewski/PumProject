���!     �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�base_estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.1.1�ub�n_estimators�K�estimator_params�(hhhhhhhhhht��	bootstrap���	oob_score���n_jobs�NhK �verbose�K �
warm_start��hN�max_samples�NhhhNhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h)�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�battery_power��blue��clock_speed��dual_sim��fc��four_g��
int_memory��n_cores��pc��ram��	talk_time��three_g��touch_screen��wifi�et�b�n_features_in_�K�
n_outputs_�K�classes_�h(h+K ��h-��R�(KK��h2�i8�����R�(K�<�NNNJ����J����K t�b�C                              �t�b�
n_classes_�K�base_estimator_�h	�estimators_�]�(h)��}�(hhhhhNhKhKhG        hh$hNhJ�
hG        hNhG        hHKhIKhJh(h+K ��h-��R�(KK��h2�f8�����R�(KhRNNNJ����J����K t�b�C               �?       @      @�t�bhVh&�scalar���hQC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh(h+K ��h-��R�(KK��hQ�C       �t�bK��R�}�(hK�
node_count�M7�nodes�h(h+K ��h-��R�(KM7��h2�V56�����R�(Kh6N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h�hQK ��h�hQK��h�hQK��h�hbK��h�hbK ��h�hQK(��h�hbK0��uK8KKt�b�B�               
            �3@ףp=
��?�            �@                          @�m�����?�           ܗ@       b                    �?ޓ�i���?P           H�@       ]                    @�
J��L�?h             g@              
             !@��5��?_             e@              	            ��@a�ʤC��?'            �Q@              
             @z�G�z�?             9@                           .�@�LQ�1	�?             7@	       
       	            h�@�C��2(�?             6@������������������������       �                     1@                           �?���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                           @\1�K36�?             G@              	            �@�8��8��?             8@                           l�@      �?              @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @                           @�@      �?	             0@������������������������       �                     �?������������������������       �                     .@                           ,�@���7�?             6@������������������������       �                     1@                           r�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @       $                    -@���C��?8            �X@        !       
             /@@4և���?             ,@������������������������       �                     &@"       #                    &@�q�q�?             @������������������������       �                     �?������������������������       �                      @%       P       
            �0@߀2q�{�?2             U@&       /                    �?��K��?'            �M@'       (       	            ؐ@�y5�h�?             >@������������������������       �                      @)       .       	            �@ˠT�x�?             6@*       +                    �?��S�ۿ?             .@������������������������       �                     &@,       -                    ��@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @0       ;                    �?ܷ��?��?             =@1       :       
             -@�(ݾ�z�?             *@2       3                    @�n���?             "@������������������������       �                     @4       9                    �?�q�q�?             @5       8                    �?z�G�z�?             @6       7                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                     @<       M                    �?      �?             0@=       B       
             '@�������?             (@>       ?                 `ff�?      �?             @������������������������       �                     �?@       A                 @33�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?C       F       
             )@�8��8��?             @D       E                   �?      �?              @������������������������       �                     �?������������������������       �                     �?G       J                    �?      �?             @H       I                    �@      �?              @������������������������       �                     �?������������������������       �                     �?K       L       
             +@      �?              @������������������������       �                     �?������������������������       �                     �?N       O       	            :�@      �?             @������������������������       �                     @������������������������       �                     �?Q       V                    x�@��ׁsF�?             9@R       S                    @h/�����?             "@������������������������       �                     @T       U                   �F@z�G�z�?             @������������������������       �                     @������������������������       �                     �?W       \                    B@     ��?             0@X       [                    <@:/����?             @Y       Z       	            ��@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     "@^       _       	            �@�.�?��?	             .@������������������������       �                     "@`       a                   @K@r�q��?             @������������������������       �                     @������������������������       �                     �?c       �       
             @b�x���?�           ��@d       }                    ,@�.�s�?             C@e       p                    �@��7S��?            �@@f       i                    �?������?             .@g       h                 hff�?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?j       o                    @���Q��?             @k       n                    �?�q�q�?             @l       m                    J@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @q       t                    �?2�tk~X�?             2@r       s                 033�?      �?              @������������������������       �                     @������������������������       �                      @u       z       	            z�@���(\��?	             $@v       w                    @؇���X�?             @������������������������       �                     @x       y                   �H@      �?              @������������������������       �                     �?������������������������       �                     �?{       |       	            ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @~       �                    �?{�G�z�?             @       �       	            Z�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�             
             #@������?�           X�@�       �                   @F@$Uކ�?�            `s@�       �                    ~�@�K�_�?�            �l@�       �                    �?���|�?P             _@�       �       	            �@=[y���?             1@�       �                    �?r�q��?
             (@�       �                    �?      �?              @�       �                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                 pff@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                 ����?��� �?D            �Z@�       �                    �?t�E]t�?             &@�       �       	            1�@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                    �?{�G�z�?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �       	            :�@r�q��?=             X@�       �                    �@P���Q�?             D@������������������������       �                    �@@�       �                    @����X�?             @�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �       	            ��@>4և���?%             L@�       �       	            �@	���ĳ�?             >@�       �                   �0@z�G�z�?	             $@�       �                    ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �?H�z�G�?             4@�       �       
             @      �?              @�       �                    !@z�G�z�?             @������������������������       �                     @�       �                 `ff@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       
             @�8��8��?             (@������������������������       �                     $@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 pff@ ��WV�?             :@������������������������       �                     9@������������������������       �                     �?�       �       	            �@�A�A�?B            @Z@�       �                    @��Q��?#             I@�       �       	            ơ@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                 033�?�2�@�4�?            �D@�       �                    @���ʻ��?             1@������������������������       �                     �?�       �                   �:@     ��?             0@������������������������       �                     $@�       �                    >@�8��8��?             @�       �       	            (�@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?�       �                    �?�������?             8@�       �       	            t�@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?h/�����?             2@�       �                    �?�z�G��?             $@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	            ?�@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �       	            (�@      �?              @������������������������       �                     �?�       �                 033�?؇���X�?             @�       �                   @B@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                    �K@�       �                 ����?�c 6���?7            @T@�       �       	            ��@������?             5@�       �                     @$�q-�?             *@������������������������       �                     �?������������������������       �                     (@�       �                    @      �?              @�       �                    �?      �?             @������������������������       �                      @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @      �?             @������������������������       �                      @�       �                   �L@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?^n����?)             N@�       �                    `�@�q�q�?             8@������������������������       �                     @�       �                    @ )O��?             2@�       �                    �?      �?              @������������������������       �                      @�       �       	            ��@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �       	            ��@ףp=
��?             $@�       �                    &@      �?              @�       �                    @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�             	            ��@�������?             B@�             	            f�@      �?             8@                          @      �?             (@������������������������       �                     "@������������������������       �                     @                         @      �?             (@������������������������       �                     @            	            Q�@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �        
             (@	      �                   �?8�.��?           Py@
                         #@�>|���?�            `i@                         @x�5?,R�?             B@                         @0��b�/�?
             .@                         d�@����X�?             @������������������������       �                     �?                         0�@r�q��?             @������������������������       �                     @            
             /@�q�q�?             @������������������������       �                     �?������������������������       �                      @            	            ��@      �?              @������������������������       �                     @                         @      �?             @������������������������       �                      @������������������������       �                      @            	            �@���N8�?             5@������������������������       �                     �?������������������������       �                     4@      K                   �?ZIY~��?o            �d@      J      	            w�@Ztjط}�?1            @R@      G                   ��@�FX�i��?$             M@      F                  �J@9��8���?             H@       5      
             +@�%�܅�?            �D@!      ,                   ��@VUUUUU�?             2@"      #                033�?��E���?             "@������������������������       �                     �?$      '                   @      �?              @%      &                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @(      +                   �?z�G�z�?             @)      *                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @-      4                   �?|	�%���?             "@.      /                   �?
ףp=
�?             @������������������������       �                      @0      1                   �?VUUUUU�?             @������������������������       �                     �?2      3                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @6      ;      	            Γ@�nkK�?             7@7      8      	            l�@"pc�
�?             &@������������������������       �                     @9      :                  @@@���Q��?             @������������������������       �                      @������������������������       �                     @<      C                   �?�q�q�?             (@=      >      
             /@      �?              @������������������������       �                     @?      @                    @���Q��?             @������������������������       �                      @A      B      	            ݥ@�q�q�?             @������������������������       �                      @������������������������       �                     �?D      E      
             1@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @H      I                  @E@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     .@L      Y                   @���}!�?>            �W@M      V      	            Z�@�X���?             6@N      O                   &@H�z�G�?
             $@������������������������       �                     �?P      Q                `ff�?�q�q�?	             "@������������������������       �                     @R      U                   �?      �?             @S      T                  �3@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @W      X                   @�8��8��?             (@������������������������       �                     �?������������������������       �                     &@Z      �                   J�@�a�2�t�?/             R@[      z                   �?���{���?+            �P@\      o                033�?     P�?             @@]      b                   @����p9�?             3@^      a                   �?���Q��?             @_      `                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @c      l                033�?���>4��?             ,@d      i      	            ѡ@b���i��?	             &@e      h                ����?�$I�$I�?             @f      g                   @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @j      k                   �?      �?             @������������������������       �                     �?������������������������       �                     @m      n                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?p      q      
             +@޾�z�<�?             *@������������������������       �                     @r      u                   @X�<ݚ�?             "@s      t                   @      �?              @������������������������       �                     �?������������������������       �                     �?v      w                   �?؇���X�?             @������������������������       �                     @x      y                   @      �?             @������������������������       �                     @������������������������       �                     �?{      �                   �?�_��*�?            �A@|      �                033�?�[��"e�?	             2@}      ~                   @������?             .@������������������������       �                      @      �                   �@և���X�?             @������������������������       �                     @�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?�      �                   :�@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   @�������?             1@�      �                   ��@$I�$I��?             ,@������������������������       �                      @�      �                  @A@      �?             (@������������������������       �                     @�      �                   '@      �?             @������������������������       �                     @������������������������       �                     @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   '@z�G�z�?             @�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   @~����?�            @i@�      �      
             )@Ӟ����?D            �Z@�      �                   -@�3�R��?             C@�      �                   &@�[���q�?             ?@�      �      	            ��@�8��8��?             8@�      �                   �?���k���?             &@������������������������       �                      @�      �                   ��@�<ݚ�?             "@������������������������       �                     @�      �                   �?      �?             @������������������������       �                      @������������������������       �                      @�      �      	            ��@$�q-�?	             *@������������������������       �                     $@�      �      
             %@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?����X�?             @�      �      	            Ο@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�      �      	            8�@����X�?             @������������������������       �                     @������������������������       �                      @�      �      	            �@7R��h`�?+            @Q@�      �                   N�@:ɨ��?            �@@�      �      
             /@�C��2(�?             6@������������������������       �                     *@�      �                   �@�<ݚ�?	             "@������������������������       �                     @�      �                   9@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?���!pc�?             &@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �      
             -@      �?              @������������������������       �                     �?������������������������       �                     @�      �                   @�"e����?             B@�      �                   @V��6���?
             1@������������������������       �                     @�      �      	            V�@���k���?             &@�      �                   �?�<ݚ�?             "@�      �                   �?���Q��?             @������������������������       �                      @�      �                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                   �?D�n�3�?             3@������������������������       �                     @�      �                   n�@�n_Y�K�?             *@������������������������       �                      @������������������������       �                     @�      �      	            ��@����p9�?=            �W@�      �                   �@ףp=
��?#             I@�      �      
             &@�X�C�?             <@�      �                    @���Q��?             @�      �                   @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�      �                   +@I�O���?             7@�      �                   0�@      �?	             0@������������������������       �                      @�      �                ����?      �?              @�      �      
             +@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �      	            ��@������?             @������������������������       �                     @�      �                   >@      �?             @������������������������       �                     @������������������������       �                     �?�      �                pff�?�X���?             6@�      �      	            ��@���k���?	             &@�      �                   �?      �?             @�      �                   @�q�q�?             @�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �?"pc�
�?
             &@�      �      	            b�@����X�?             @������������������������       �                     @������������������������       �                      @�      �                   �?      �?             @�      �                   �?�q�q�?             @������������������������       �                     �?�      �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�                         B@�<ݚ�?            �F@�            	            ��@���7�?             6@�                          �?z�G�z�?             @�      �      
             .@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        	             1@                        �D@�û��|�?             7@������������������������       �                     @                         �?�d�����?             3@                         �?X�<ݚ�?             "@������������������������       �                     @                         �?z�G�z�?             @	      
                   @�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @            
             '@ףp=
�?             $@                        �M@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @      _      	            4�@�5IYp��?o           p�@      ^                  �O@�1�=B��?�            @o@      M                033�?W��dִ�?�            `n@      (                   ��@��_?WQ�?c            �c@                         @�����?$            �L@������������������������       �                     @                         @Ȩ�I��?#            �J@                         �?p�ݯ��?             3@������������������������       �                     @            	            ��@z�G�z�?	             .@������������������������       �                     (@������������������������       �                     @      '                   M@H�V�e��?             A@                          -@     ��?             @@������������������������       �                     "@!      &      	            ��@��<b���?             7@"      #                   @�}�+r��?             3@������������������������       �        	             .@$      %      
             +@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @)      6      	            r�@�BD`�z�??            @Y@*      1                   ��@��k=.��?            �G@+      0                   @�8��8��?             B@,      -                   �?�q�q�?             "@������������������������       �                     @.      /                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ;@2      3      	            �}@�eP*L��?             &@������������������������       �                      @4      5                   �?�q�q�?             "@������������������������       �                     @������������������������       �                     @7      F                   )@H�ՠ&��?#             K@8      A                   @����X�?             5@9      :                  @@@�eP*L��?             &@������������������������       �                     �?;      <                   x�@���Q��?             $@������������������������       �                     @=      >      	            R�@�q�q�?             @������������������������       �                     @?      @                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @B      C                   @ףp=
�?             $@������������������������       �                     @D      E                   �?      �?             @������������������������       �                     @������������������������       �                     �?G      H                   �?Pa�	�?            �@@������������������������       �                     2@I      L                  �0@��S�ۿ?
             .@J      K                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@N      W                  �2@vQ-	���?3            @U@O      P      	            ��@     �?(             P@������������������������       �                     G@Q      R                   �@b�2�tk�?             2@������������������������       �                     @S      T                   %@$�q-�?	             *@������������������������       �                     &@U      V      	            J�@      �?              @������������������������       �                     �?������������������������       �                     �?X      Y                   t�@����X�?             5@������������������������       �                     @Z      [                   �?      �?             0@������������������������       �                     &@\      ]                  �J@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @`      �                `ff@#)/5;A�?�            @u@a      �                  �6@����
�?�            �q@b      �                   z�@;����?G             [@c      �      	            ��@tv?z���?<            �V@d      i                ����?�~E�0��?1             S@e      f                   �?b�2�tk�?             2@������������������������       �                      @g      h      
             !@�z�G��?             $@������������������������       �                     @������������������������       �                     @j      q                   �?���d�?%             M@k      l      	            �@������?             @������������������������       �                     @m      p                   @      �?             @n      o                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @r      u      
             @L紂P�?             �I@s      t                   h�@և���X�?             @������������������������       �                     @������������������������       �                     @v      }      
             !@t��ճC�?             F@w      x                `ff�?z�G�z�?
             $@������������������������       �                     @y      |                   @�q�q�?             @z      {      	            p�@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @~                         @г�wY;�?             A@������������������������       �                    �@@������������������������       �                     �?�      �      
             #@؇���X�?             ,@�      �                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�      �                   ֝@X�<ݚ�?             2@�      �                   @���!pc�?             &@������������������������       �                      @������������������������       �                     @�      �                   �?����X�?             @������������������������       �                     �?�      �                ����?r�q��?             @������������������������       �                     �?������������������������       �                     @�      �                   �@��K���?q            `f@�      �                   �?��8��8�?             (@�      �      
             "@���Q��?             @������������������������       �                      @�      �                  �:@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �      	            ��@��		�?j            �d@�      �                   !@�#N�?A            �Y@�      �                  �;@�<ݚ�?'            �O@�      �                   �?      �?             @�      �      	            ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �                `ff�?6N���?$            �M@�      �                   �?�g���e�?	             &@������������������������       �                     @�      �                   @������?             @������������������������       �                     @�      �                   �?      �?             @������������������������       �                      @�      �                   @�@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                `ff @r�qG�?             H@�      �                  �3@T���N@�?             9@�      �                   �? �q�q�?             8@������������������������       �                     4@�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   !@��<b���?             7@�      �                   @�q�q�?             @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �      
             @�IєX�?             1@�      �                  �J@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@�      �                  �2@p=
ףp�?             D@�      �                033@     ��?             @@�      �                   b�@�-Z�?             =@�      �      
             @�z�G��?             4@������������������������       �                     @�      �                   @@��
ц��?
             *@������������������������       �                     @�      �                   �?      �?              @�      �                   @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�      �      
              @�����H�?             "@������������������������       �                     �?������������������������       �                      @�      �                   @�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?      �?              @������������������������       �                      @�      �                   @�q�q�?             @������������������������       �                     @������������������������       �                      @�      �                   �?      �?)             P@�      �      
             &@�>4և��?             <@�      �                ����?�����?             5@�      �      
             @���Q��?             @������������������������       �                      @�      �                   @�q�q�?             @������������������������       �                     �?�      �      	            ʫ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             0@�      �      	            ��@և���X�?             @������������������������       �                      @�      �                  �K@z�G�z�?             @�      �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   @�8��8��?             B@�      �                   �?@�0�!��?             1@�      �                  �J@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                  @@@�8��8��?	             (@�      �                   1@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �        	             3@�      �      
             @ZhZ�-�?            �J@�      �                   l�@�����H�?             "@������������������������       �                     �?������������������������       �                      @�                         )@5_�g���?             F@�            	            i�@��	"P7�?             C@�                        �3@lxz�,C�?             9@�      �      
             -@      �?             8@�      �      
             (@�S����?
             3@������������������������       �                     @�      �                   �?�θ�?             *@�      �                   /@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�                          @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@������������������������       �                     @                         ?@.*��\�?/            @R@                         �?yA+��?            �C@      
                   �?=[y���?             1@      	                   @      �?              @������������������������       �                     @������������������������       �                     @                         �?X�<ݚ�?             "@������������������������       �                     @                         Č@�q�q�?             @������������������������       �                      @������������������������       �                     �?                         +@��#��Z�?             6@                         @     ��?
             0@            	            "�@����S�?	             ,@                         d�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@������������������������       �                      @            	            ǣ@      �?             @������������������������       �                     @������������������������       �                     @      &                   �?>z��.k�?             A@                         �?���(\��?             $@������������������������       �                     @                         �?�q�q�?             @������������������������       �                     �?       #                    @{�G�z�?             @!      "                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @$      %                   �@      �?              @������������������������       �                     �?������������������������       �                     �?'      .                  �J@�q�q�?             8@(      -      	            0�@x�5?,�?             "@)      *                   �?r�q��?             @������������������������       �                     @+      ,                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @/      4      	            ��@*;L]n�?             .@0      3                   ,@�C��2(�?             &@1      2      	            t�@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @5      6                   �?      �?             @������������������������       �                      @������������������������       �                      @�t�b�values�h(h+K ��h-��R�(KM7KK��hb�B�f       x@     �w@     �z@     Py@     pw@     v@     @z@     �w@      n@     �h@      n@     0p@     �P@      =@     �F@     �E@      M@      =@      D@      E@      4@      @      <@      0@      4@      @                      4@      @                      4@       @                      1@                              @       @                      @                                       @                              �?                               @                               @      <@      0@               @      @      .@               @      @                       @      �?                       @                                      �?                              @                              �?      .@                      �?                                      .@                      5@      �?                      1@                              @      �?                              �?                      @              C@      6@      (@      :@      *@                      �?      &@                               @                      �?                              �?       @                              9@      6@      (@      9@      2@      6@      @      *@      "@      ,@              @       @                              �?      ,@              @      �?      ,@                              &@                      �?      @                              @                      �?                                                      @      "@       @      @      @      @      @      @       @      @      @               @      @                                      @               @              @              �?               @              �?                              �?               @                               @                                              �?                      @              @      @       @      @      @      @      �?      @      �?      �?              @              �?                      �?                      @                              @      �?                               @      @      �?                      �?      �?                              �?                      �?                       @       @                      �?      �?                              �?                      �?                              �?      �?                      �?                                      �?                      @              �?              @                                              �?              @              @      (@      @              @      �?                      @              @                      �?      @                                                      �?      @               @      &@      @               @       @                       @       @                       @                                       @      @                                                      "@      "@              @      �?      "@                                              @      �?                      @                                      �?     �e@     �d@     �h@      k@      @      $@      2@      @      @       @      2@       @      @              &@              �?              "@                              "@              �?                              @               @              �?               @              �?              �?              �?                                              �?                              �?               @                              �?       @      @       @               @      @                              @                       @                      �?      @      �?       @      �?      @                              @                      �?      �?                              �?                      �?                                              �?       @                      �?                                       @      �?       @               @      �?       @                      �?                                       @                                               @      e@     �c@     @f@     �j@     �R@      P@      O@     @[@      J@      E@     �F@     �V@     �E@      8@      8@     �@@       @      "@      �?      @       @      "@      �?               @      @      �?                      @      �?                      @                                      �?               @      �?                       @                                      �?                              @                                              @     �D@      .@      7@      <@      �?      �?      @       @      �?              @              �?                                              @                      �?       @       @              �?                                       @       @                               @                       @              D@      ,@      0@      :@      C@       @                     �@@                              @       @                      �?       @                      �?                                       @                      @                               @      (@      0@      :@       @      (@      .@      �?       @       @                       @      �?                       @                                      �?                              @                              @      .@      �?              @      @                      �?      @                              @                      �?      �?                              �?                      �?                              @                                      &@      �?                      $@                              �?      �?                              �?                      �?                              �?      9@                              9@                      �?              "@      2@      5@     �L@      "@      2@      5@       @              @       @                      @                                       @              "@      &@      3@       @      @      �?      (@      �?              �?                      @              (@      �?                      $@              @               @      �?      @               @              @                                               @                                      �?      @      $@      @      �?      @      �?                      @                                      �?                      �?      "@      @      �?              @      @                       @      �?                       @                                      �?                      �?      @                      �?                                      @              �?      @              �?      �?                                      @              �?              �?              �?                              �?              �?                              @                                             �K@      7@      6@      1@      3@      (@      @      @      @      (@      �?                              �?                      (@                                       @      @      @              �?      @                               @                      �?      �?                              �?                      �?                              �?              @                               @              �?              �?              �?                                              �?      &@      3@      ,@      0@       @      @      &@      @                      @               @      @      @      @       @      @               @       @                                      @               @              @                                               @              @      @       @              @      @                      �?      @                              @                      �?                               @                                               @      "@      (@      @      (@      "@      (@      @              "@      @                      "@                                      @                              "@      @                      @                              @      @                      @                                      @                                      (@     @W@     @W@      ]@     �Y@      H@      F@     �Q@     �D@      @       @      9@       @      @       @      @       @       @              @              �?                              �?              @                              @              �?               @              �?                                               @              @       @               @      @                                       @               @               @                                               @      �?              4@              �?                                              4@             �D@      E@     �F@     �C@      2@      9@      (@      2@      2@      9@      (@      @      2@      0@      (@       @      &@      0@      (@       @       @      @       @       @      �?      @       @      �?                              �?      �?      @       @                      �?       @                      �?                                       @              �?      @                      �?       @                               @                      �?                                       @                      �?      �?      @      �?      �?      �?       @      �?                       @              �?      �?              �?                              �?      �?      �?                      �?                                      �?                                      @              "@      $@      @              "@       @                      @                              @       @                               @                      @                                       @      @                      @      @                      @                               @      @                               @                       @      �?                       @                                      �?                      @      �?                              �?                      @                      @                                      "@              �?              "@                                              �?                              .@      7@      1@     �@@      5@      @      @       @      &@      @      @      �?                              �?              @      @                      @                              @      @                      @      �?                              �?                      @                                       @                                      �?      &@                      �?                                      &@      1@      ,@      ?@      $@      1@      $@      ?@      "@      @       @      ,@      @      @      @      @      @              @               @              �?               @                               @              �?                               @                      @      @      @      @      �?      @      @      @      �?      @       @              �?               @              �?                                               @                      @                                      �?      @                      �?                                      @       @              �?               @                                              �?               @      �?      $@                              @               @      �?      @              �?      �?                              �?                      �?                              �?              @                              @              �?              @                              @              �?                              (@       @      1@      @      @              &@      �?      @              &@                               @              @              @              @                              �?              @                              @              �?                               @                      �?                              �?       @                              @       @      @      @      @              @      @                       @              @              @      @      @                                              @      @                      @                                      @               @      �?                              �?                       @                              @              �?              �?              �?                              �?              �?                              @                     �F@     �H@      G@      O@      >@      8@      :@      ;@      @      (@      @      ,@       @      (@      @      (@       @      @      @      (@       @      @       @               @                                      @       @                      @                               @       @                               @                       @                                      �?      (@                              $@                      �?       @                      �?                                       @              @       @                      @       @                      @                                       @                       @                      @                       @      @                                                       @      7@      (@      5@      *@      7@      $@                      4@       @                      *@                              @       @                      @                              �?       @                      �?                                       @                      @       @                       @      �?                              �?                       @                              �?      @                      �?                                      @                               @      5@      *@               @      *@       @                      @                       @      @       @               @      @                       @      @                               @                       @      �?                       @                                      �?                              @                                       @                       @      &@                              @                       @      @                       @                                      @      .@      9@      4@     �A@      .@      9@      $@              @      4@      �?              @       @                      �?       @                      �?                                       @                       @                              @      2@      �?              �?      .@                               @                      �?      @                      �?       @                               @                      �?                                      @                      @      @      �?              @                                      @      �?                      @                                      �?               @      @      "@               @       @      @               @       @                      �?       @                      �?      �?                      �?                                      �?                              �?                      �?                                              @              @      @       @              @       @                      @                                       @                      �?      �?       @              �?               @                              �?              �?              �?              �?                                              �?                      �?                                      $@     �A@                      �?      5@                      �?      @                      �?      �?                      �?                                      �?                              @                              1@                      "@      ,@                      @                              @      ,@                      @      @                              @                      @      �?                       @      �?                       @                                      �?                       @                              �?      "@                      �?       @                      �?                                       @                              @     �`@     �c@     `f@      ^@     �`@      [@       @             �`@     @Y@       @             @S@     �R@      @             �C@      2@                              @                     �C@      ,@                      (@      @                              @                      (@      @                      (@                                      @                      ;@      @                      ;@      @                      "@                              2@      @                      2@      �?                      .@                              @      �?                      @                                      �?                              @                               @                      C@      L@      @              C@      "@                     �@@      @                      @      @                      @                              �?      @                              @                      �?                              ;@                              @      @                       @                              @      @                      @                                      @                             �G@      @                      .@      @                      @      @                              �?                      @      @                      @                               @      @                              @                       @      �?                              �?                       @                              "@      �?                      @                              @      �?                      @                                      �?                      @@      �?                      2@                              ,@      �?                      @      �?                      @                                      �?                      &@                     �L@      ;@      �?             �I@      (@      �?              G@                              @      (@      �?              @                                      (@      �?                      &@                              �?      �?                      �?                                      �?              @      .@                      @                              �?      .@                              &@                      �?      @                              @                      �?                                      @                             �H@     `e@      ^@             �F@      c@     @V@              1@      Q@      7@              1@      N@      *@              1@      M@      �?              @      &@                               @                      @      @                              @                      @                              $@     �G@      �?              @      @      �?              @                                      @      �?                      �?      �?                              �?                      �?                               @                      @      F@                      @      @                      @                                      @                      @     �D@                       @       @                              @                       @      @                       @       @                       @                                       @                               @                      �?     �@@                             �@@                      �?                                       @      (@                       @      @                              @                       @                                       @                       @      $@                      @       @                               @                      @                              @       @                              �?                      @      �?                              �?                      @                      <@     @U@     �P@              @       @      @                       @      @                               @                       @      �?                              �?                       @                      @                              5@     �T@     �O@              5@     �R@      @              "@      I@      @                       @       @                      �?       @                      �?                                       @                      �?                      "@      H@       @              @      @      �?                      @                      @      @      �?                      @                      @              �?               @                              �?              �?              �?                                              �?              @     �D@      �?              �?      7@      �?                      7@      �?                      4@                              @      �?                              �?                      @                      �?                              @      2@                      @       @                      �?       @                      �?                                       @                      @                              �?      0@                      �?       @                      �?                                       @                              ,@                      (@      9@      @               @      7@      �?              @      6@      �?              @      ,@                              @                      @      @                              @                      @       @                       @       @                       @                                       @                      @                                       @      �?                              �?                       @                       @      �?                              �?                       @                              @       @       @                       @                      @               @              @                                               @                       @      L@                      @      7@                       @      3@                       @      @                               @                       @      �?                      �?                              �?      �?                      �?                                      �?                              0@                      @      @                       @                              �?      @                      �?      �?                              �?                      �?                                      @                      @     �@@                      @      ,@                       @      @                              @                       @                              �?      &@                      �?       @                               @                      �?                                      "@                              3@              @      2@      ?@              �?               @              �?                                               @              @      2@      7@              @      2@      1@              @      2@      @              @      2@      @                      0@      @                      @                              $@      @                      @      @                              @                      @                              @                      @       @                      @                                       @                                      �?                              *@                              @      $@      ;@      $@      :@      @      .@      �?      4@       @      "@      �?      @              @              @              @                                              @       @      @      �?                      @                       @              �?               @                                              �?              �?      @              .@      �?      @              (@      �?      �?              (@      �?      �?                      �?                                      �?                                              (@               @                              @              @              @                                              @      @      (@      "@      @      @      �?       @      �?      @                               @      �?       @      �?                              �?       @      �?       @              �?               @              �?                                               @              �?      �?                      �?                                      �?                      �?      &@      @      @              �?      @      @              �?      @                              @                      �?      �?                      �?                                      �?                                      @      �?      $@       @       @      �?      $@                      �?      @                      �?                                      @                              @                                       @       @                               @                       @        �t�bub��r     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJ/��hG        hNhG        hHKhIKhJh(h+K ��h-��R�(KK��hb�C               �?       @      @�t�bhVhghQC       ���R�hkKhlhoKh(h+K ��h-��R�(KK��hQ�C       �t�bK��R�}�(hKhyMChzh(h+K ��h-��R�(KMC��h��B�~         H      	            R�@���&��?�            �@       �                    d�@4C�?�?�           ��@       �                    �?H�uh)��?�           ��@       '                    �?Yv�3Q�?�            �t@       
                 ����?��wvJ�?3            �V@                           �?�IєX�?             1@������������������������       �                     (@       	                    �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?                           H@rH\O���?+            @R@                           �?d}h���?              L@                           @�q�q�?             (@              	            p�@���Q��?             @������������������������       �                      @������������������������       �                     @              	            r�@؇���X�?             @������������������������       �                     �?������������������������       �                     @                           ��@�C��2(�?             F@                           x�@z�G�z�?	             .@������������������������       �                     $@                           @���Q��?             @                            @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @              	            �@XB���?             =@������������������������       �                     <@������������������������       �                     �?       $                    @.k��\�?             1@        #                 ����?$�q-�?             *@!       "       
             $@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     "@%       &                    @      �?             @������������������������       �                     @������������������������       �                     �?(       q                    @�Gӹ�?�            �n@)       T                    @��J�-�?p            �f@*       A                    �?��'��
�?E            �[@+       >                    .@S)Vr!��?%            @P@,       -                    @NI��&�?"             M@������������������������       �                     @.       9       	            B�@n�7{P��?            �K@/       0       	            ��@�}�+r��?             C@������������������������       �                     ;@1       8                    �?"pc�
�?             &@2       3                    �?����X�?             @������������������������       �                     @4       7                    @�q�q�?             @5       6                    ,@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @:       =                    �?@�0�!��?
             1@;       <                   �3@�q�q�?             "@������������������������       �                     @������������������������       �                     @������������������������       �                      @?       @       
             $@����X�?             @������������������������       �                     @������������������������       �                      @B       C       	            ��@�nkK�?              G@������������������������       �        
             .@D       Q                 ��� @�?Q�f?�?             ?@E       F                    $@      �?             8@������������������������       �                     @G       H                    �?؇���X�?             5@������������������������       �                     &@I       J                    )@�z�G��?             $@������������������������       �                      @K       L                    .@      �?              @������������������������       �                     �?M       P                   �:@����X�?             @N       O                    v�@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                      @R       S                    ��@����X�?             @������������������������       �                      @������������������������       �                     @U       ^                    +@F��ӭ��?+             R@V       ]                    ��@�z�G��?             4@W       X                    @      �?             (@������������������������       �                     @Y       \       
             !@      �?              @Z       [                    @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @_       b       
             @�E��
��?             J@`       a       	             �@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@c       f                    @      �?             D@d       e       	            ,�@և���X�?	             ,@������������������������       �                      @������������������������       �                     @g       h                    �?8�Z$���?             :@������������������������       �                     @i       p       
            �3@���y4F�?
             3@j       o                    �@r�q��?	             2@k       n                    t�@���Q��?             @l       m       	            j�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                     �?r       w       
             !@�jTM��?$            �N@s       v       
             @Pa�	�?            �@@t       u                 033@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ;@x       �                 pff@      �?             <@y       |                 `ff�?�q�q�?             5@z       {                    '@      �?             @������������������������       �                     @������������������������       �                     �?}       �                   @N@������?             1@~                           �?�r����?
             .@������������������������       �                      @�       �       	            ~�@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �       	            ��@I�9v�'�?�            @t@�       �                   @F@J� ��w�?s             g@�       �       	            r�@�L�w��?V            �a@�       �                    �@���F6��?<            �X@�       �                    �?����ȫ�?2            �T@�       �                    @r�q��?             @�       �                    -@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �        -             S@�       �                    ��@ҳ�wY;�?
             1@�       �                   �C@z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    �?r�q��?             (@������������������������       �                     $@������������������������       �                      @�       �                    @D^��#��?            �D@�       �                   �;@      �?             8@�       �                    �?�q�q�?             2@�       �                 (33�?����X�?             @�       �                 ����?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?�C��2(�?             &@������������������������       �                      @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �                    �@������?             1@������������������������       �        	             *@������������������������       �                     @�       �       	            ��@`���i��?             F@������������������������       �                     D@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �       
            �3@�ǫz��?Z            �a@�       �                   �I@��a!�z�?U            �`@�       �                    #@,ҭb���?H            @\@�       �                    �?4;�Wp��?=            @X@�       �                    �@�bC�B��?"            �H@�       �                    �?���Q��?             @������������������������       �                      @�       �                    ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                 pff�?N�zv�?             F@�       �       
            �1@T���N@�?             9@�       �                    @���7�?             6@�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@�       �       	            ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @B+K&:~�?             3@�       �       
             &@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    !@H�7�&��?             .@�       �                    @؇���X�?
             ,@������������������������       �                      @������������������������       �        	             (@������������������������       �                     �?�       �                    �?@��8��?             H@�       �                    @��S�ۿ?	             .@�       �                    �?؇���X�?             @������������������������       �                     @�       �       
             '@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                    �@@�       �                    `�@      �?             0@�       �                    �?r�q��?	             (@�       �                    6@����X�?             @������������������������       �                     @�       �                    ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �                   �J@R��Xp�?             3@������������������������       �                     @�       �                 033�?������?             .@�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @�       �       	            b�@�C��2(�?	             &@�       �                   �L@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�       �                   @M@      �?              @������������������������       �                     @�       �                    ̎@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?j�n`��?j            �d@�       �                    �?�[��"e�?             2@�       �                    �?��8��8�?             (@�       �                    @X�<ݚ�?             "@�       �                    B�@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�                          6@Y�V��7�?b            �b@�                          @N<+	��?&             N@�       �       
             @���n(T�?            �@@�       �       	            ��@�q�q�?             (@������������������������       �                     @������������������������       �                     @�                          @�E�_���?             5@�                          &@B{	�%��?             "@                          +@      �?              @������������������������       �                     @                         @      �?             @������������������������       �                      @                         �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@	            
             /@;����?             ;@
                         .@�lO���?
             3@            	            ؏@      �?             (@������������������������       �                     @������������������������       �                     @                         �?����X�?             @������������������������       �                     �?                         �?r�q��?             @������������������������       �                     @������������������������       �                     �?                         �?      �?              @������������������������       �                      @������������������������       �                     @      E                   @&ޏ���?<             V@      ,                   @
�Sy'�?8             U@      #                   @hE#߼�?            �F@      "                   �?@�0�!��?             A@                         @ҳ�wY;�?             1@������������������������       �                      @      !      
            �1@�q�q�?             "@                         �?؇���X�?             @������������������������       �                     @                          F@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     1@$      %      	            X�@��ˠ�?             &@������������������������       �                     @&      '                   �?      �?              @������������������������       �                      @(      +                  @D@r�q��?             @)      *      
            �1@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @-      .      
             @�V��B�?            �C@������������������������       �                     @/      >                ����?f�t���?             A@0      7                   ��@V����?             6@1      4                   @{�G�z�?             $@2      3                   ��@���Q��?             @������������������������       �                     @������������������������       �                      @5      6                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @8      9                   �?�������?	             (@������������������������       �                     @:      ;                ����?�Q����?             @������������������������       �                     @<      =                   �?      �?              @������������������������       �                     �?������������������������       �                     �??      @                   '@r�q��?	             (@������������������������       �                      @A      D                   �?      �?             @B      C      
             &@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @F      G                   ��@      �?             @������������������������       �                     �?������������������������       �                     @I      �      	            ��@��ΑQ��?�           @�@J      �                   Ԕ@x 5?6>�?�            `w@K      �                   '@��I�?�            �l@L      i      	            �@ji_}a�?�            �j@M      b                   @8tM���?#            �L@N      S      	            
�@�'���{�?             G@O      R                   x�@      �?
             0@P      Q                   �?����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     "@T      ]                  �K@z5�h$�?             >@U      \                   �?D%��N��?             7@V      [      	            �@H�z�G�?             $@W      Z                   �?�8��8��?             @X      Y                ����?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     *@^      a                   @����X�?             @_      `                   �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?c      h      
             /@���|���?             &@d      g                   ,@�<ݚ�?             "@e      f                   @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @j      �      
             /@�#}w���?b            �c@k      ~                   @�#3����?J             ]@l      w      	            ͤ@,�T�6�?A             Z@m      r                   ��@R���Q�?             D@n      o                   @����X�?             @������������������������       �                     @p      q      	            Q�@�q�q�?             @������������������������       �                     �?������������������������       �                      @s      v                   �?Pa�	�?            �@@t      u                   @r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ;@x      }                   �?     ��?&             P@y      z      
             %@$�q-�?             *@������������������������       �                     $@{      |      	            E�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                    �I@      �      
             "@�q�q�?	             (@�      �                  �A@r�q��?             @������������������������       �                     @�      �                   H@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   0@      �?             @������������������������       �                     @������������������������       �                     @�      �                   @$6M5��?            �D@�      �                   �?ףp=
��?             $@�      �      
             2@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�      �                   �?��a�n`�?             ?@�      �                   @`2U0*��?             9@�      �                  �2@؇���X�?             @�      �      	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        	             2@�      �                   �?�q�q�?             @�      �                   �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�      �      
             @f�t���?
             1@������������������������       �                      @�      �                   -@�<ݚ�?             "@������������������������       �                      @������������������������       �                     @�      �                   ��@|�����?T            �a@�      �                   �@      �?             (@������������������������       �                     @�      �                   +@      �?              @�      �                   �?����X�?             @�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?z�G�z�?             @�      �      	            �@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?�      �                   #@���ā�?M            ``@�      �      	            �@������?@            @Z@�      �      
            �2@\���(��?-             T@�      �                ����?o%W�?'            �Q@�      �                  �G@     ��?             @@�      �                  �<@$�q-�?             :@������������������������       �        
             0@�      �      	            �@z�G�z�?             $@������������������������       �                     �?�      �                   @�����H�?             "@������������������������       �                      @������������������������       �                     �?�      �                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @�      �                   0�@��Ha���?            �C@�      �                   �?      �?              @������������������������       �                     @������������������������       �                      @�      �                   �?�g�y��?             ?@�      �      
             @؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     8@�      �                   @X�<ݚ�?             "@�      �                   �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                   �?� �	��?             9@�      �                   @؇���X�?             @������������������������       �                     @�      �                  �A@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                  @L@X�<ݚ�?             2@�      �      
             (@�q�q�?             .@�      �                   @      �?              @������������������������       �                     �?������������������������       �                     @�      �                   �?և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�      �                   !@�	j*D�?             :@�      �                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                   )@��s����?
             5@������������������������       �                      @�      �      	            
�@�KM�]�?	             3@�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     0@�                         �?�Y����?�             y@�            	            ��@��ϓ8��?w            �h@�      �                   |�@Hث3���?.            �S@�      �                   �?:�&���?            �C@�      �                   3@�q�q�?             2@������������������������       �                     @�      �                   ,@؇���X�?             ,@������������������������       �                     "@�      �                  �O@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                   �?���N8�?             5@������������������������       �                     ,@�      �                  �:@؇���X�?             @������������������������       �                     @�      �                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?�                         �?8�Z$���?            �C@�      �      	            ��@���N8�?             5@�      �                   �?؇���X�?
             ,@�      �                   @�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     @�      �                ���@և���X�?             @������������������������       �                     @                         @L@      �?             @������������������������       �                     �?������������������������       �                     @                         '@�X�<ݺ?             2@������������������������       �                     *@                         �@z�G�z�?             @������������������������       �                     �?������������������������       �                     @            
            �2@H��ԛ�?I            �]@	                        �6@�O4R���?B            �Z@
                      ����? >�֕�?            �A@                         '@�<ݚ�?             "@������������������������       �                     @                      ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     :@������������������������       �        +            �Q@                         @�θ�?             *@                         '@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @      :                   ��@�+^Ur�?y            �i@      9      	            m�@PN���?4            @V@      8                   @b�2�tk�?'             R@      7      	            ;�@�#}7��?$            �P@      ,                   �?@i��M��?"            @P@      +                   @�ՙ/�?             E@      "                   �?��S���?             >@            	            v�@      �?             (@������������������������       �                     @       !                   @���Q��?             @������������������������       �                      @������������������������       �                     @#      *                  �@@b�2�tk�?             2@$      )                   -@�q�q�?             (@%      &                   �?����X�?             @������������������������       �                     �?'      (                   �?r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     (@-      2                   �?��<b���?             7@.      1                   �?X�<ݚ�?             "@/      0                   @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @3      6                   �?@4և���?             ,@4      5      
             @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     &@������������������������       �                      @������������������������       �                     @������������������������       �                     1@;      B      	            ��@@m���?E             ]@<      =                   �?ףp=
�?             $@������������������������       �                     @>      A                   �?z�G�z�?             @?      @                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �        ?            �Z@�t�bh�h(h+K ��h-��R�(KMCKK��hb�B`H       �y@     �x@     �x@     �x@     �y@     �u@      P@             `w@     �o@      ?@             �i@     @\@      1@             �O@      :@      �?              0@      �?                      (@                              @      �?                      @                                      �?                     �G@      9@      �?              F@      (@                      @       @                      @       @                               @                      @                              �?      @                      �?                                      @                      D@      @                      (@      @                      $@                               @      @                       @      �?                              �?                       @                                       @                      <@      �?                      <@                                      �?                      @      *@      �?                      (@      �?                      @      �?                              �?                      @                              "@                      @      �?                      @                                      �?                     �a@     �U@      0@             �W@      R@      0@              M@     �B@      0@              C@      3@       @              B@      3@      @                      @                      B@      0@      @              B@       @                      ;@                              "@       @                      @       @                      @                              �?       @                      �?      �?                              �?                      �?                                      �?                      @                                      ,@      @                      @      @                              @                      @                               @                       @              @                              @               @                              4@      2@       @              .@                              @      2@       @              @      2@      @                              @              @      2@                              &@                      @      @                               @                      @      @                      �?                               @      @                       @      @                       @                                      @                               @                       @              @               @                                              @             �B@     �A@                      @      ,@                      @      @                              @                      @       @                       @       @                               @                       @                              @                                       @                      ?@      5@                      �?      &@                      �?                                      &@                      >@      $@                       @      @                       @                                      @                      6@      @                      @                              .@      @                      .@      @                       @      @                       @      �?                       @                                      �?                               @                      *@                                      �?                      G@      .@                      @@      �?                      @      �?                      @                                      �?                      ;@                              ,@      ,@                      ,@      @                      �?      @                              @                      �?                              *@      @                      *@       @                       @                              @       @                      @                                       @                               @                              @                     @e@     �a@      ,@             @c@      >@                     �[@      =@                      W@      @                     @T@      �?                      @      �?                       @      �?                              �?                       @                              @                              S@                              &@      @                      �?      @                              @                      �?                              $@       @                      $@                                       @                      3@      6@                      @      2@                      @      (@                      @       @                       @       @                       @                                       @                      @                              �?      $@                               @                      �?       @                               @                      �?                                      @                      *@      @                      *@                                      @                     �E@      �?                      D@                              @      �?                      @                                      �?                      0@     �[@      ,@              (@     �Z@      ,@               @     �W@      $@               @     @U@      @               @      C@      @              @       @                       @                              �?       @                               @                      �?                              @      B@      @              �?      7@      �?                      5@      �?                      @      �?                      @                                      �?                      2@                      �?       @                               @                      �?                              @      *@       @              @      �?                      @                                      �?                      �?      (@       @                      (@       @                               @                      (@                      �?                                     �G@      �?                      ,@      �?                      @      �?                      @                              @      �?                      @                                      �?                       @                             �@@                              $@      @                      $@       @                      @       @                      @                              �?       @                      �?                                       @                      @                                      @              @      &@      @              @                                      &@      @                      �?      @                      �?                                      @                      $@      �?                      @      �?                              �?                      @                              @                      @      @                      @                              �?      @                      �?                                      @                      D@     @W@     �@@              &@      @      �?              @      @      �?               @      @      �?              �?      @                      �?                                      @                      �?              �?                              �?              �?                              @                              @                              =@     �U@      @@              3@      @@      "@               @      8@      �?              @      @                      @                                      @                      �?      3@      �?              �?      @      �?                      @      �?                      @                              @      �?                       @                              �?      �?                      �?                                      �?              �?                                      (@                      &@       @       @              &@      @       @              @      @                      @                                      @                      @               @                              �?              @              �?              @                                              �?                       @      @                       @                                      @              $@     �K@      7@              @      K@      7@              @     �@@      "@                      <@      @                      &@      @                       @                              @      @                      �?      @                              @                      �?       @                               @                      �?                               @                              1@                      @      @      @              @                                      @      @                               @                      @      �?                      �?      �?                      �?                                      �?                      @                      @      5@      ,@                      @                      @      0@      ,@              @      ,@      @               @      @      @               @      @                              @                       @                                      �?      @                      �?                                      @              �?      $@      �?                      @                      �?      @      �?                      @                      �?              �?              �?                                              �?              �?       @      "@                               @              �?       @      �?              �?              �?                              �?              �?                                       @                      @      �?                              �?                      @                                     �I@     �t@     �x@             �I@     0p@      P@             �H@     @e@      (@             �D@     `d@      $@              =@      ;@      �?              9@      4@      �?              ,@       @                      @       @                               @                      @                              "@                              &@      2@      �?              @      0@      �?              @      @      �?               @      @      �?                      @      �?                              �?                      @                       @                              @                                      *@                      @       @                      @      �?                              �?                      @                                      �?                      @      @                       @      @                       @      @                              @                       @                                      @                       @                              (@      a@      "@              @     @Z@      @              @     @X@      �?              @      A@                      @       @                      @                              �?       @                      �?                                       @                      �?      @@                      �?      @                              @                      �?                                      ;@                             �O@      �?                      (@      �?                      $@                               @      �?                       @                                      �?                     �I@                      �?       @      @              �?      @                              @                      �?      �?                      �?                                      �?                              @      @                      @                                      @              @      ?@      @               @      @      @               @      @                              @                       @                                              @              @      <@                      �?      8@                      �?      @                      �?      �?                      �?                                      �?                              @                              2@                       @      @                       @       @                       @                                       @                               @                       @      @       @               @                                      @       @                               @                      @                       @     @V@      J@                      @      "@                              @                      @      @                       @      @                      �?      �?                              �?                      �?                              �?      @                      �?       @                      �?                                       @                               @                      �?                       @     �U@     �E@               @     �S@      9@               @     �P@      &@               @      O@      @                      :@      @                      8@       @                      0@                               @       @                              �?                       @      �?                       @                                      �?                       @      @                              @                       @                       @      B@      �?               @      @                              @                       @                                      >@      �?                      @      �?                              �?                      @                              8@                              @      @                      �?      @                              @                      �?                              @                              &@      ,@                      �?      @                              @                      �?       @                      �?                                       @                      $@       @                      $@      @                      @      �?                              �?                      @                              @      @                      @                                      @                              @                       @      2@                      @      �?                              �?                      @                              @      1@                       @                               @      1@                       @      �?                              �?                       @                                      0@                      R@     �t@                     �E@     @c@                      C@      D@                      @@      @                      (@      @                              @                      (@       @                      "@                              @       @                      @                                       @                      4@      �?                      ,@                              @      �?                      @                               @      �?                       @                                      �?                      @     �@@                      @      0@                       @      (@                       @      @                       @                                      @                              @                      @      @                              @                      @      �?                              �?                      @                              �?      1@                              *@                      �?      @                      �?                                      @                      @     �\@                       @      Z@                       @     �@@                       @      @                              @                       @      �?                              �?                       @                                      :@                             �Q@                      @      $@                      @       @                      @                                       @                               @                      =@      f@                      <@     �N@                      <@      F@                      7@      F@                      5@      F@                      0@      :@                      0@      ,@                      "@      @                      @                               @      @                       @                                      @                      @      &@                      @      @                       @      @                      �?                              �?      @                      �?                                      @                      @                                      @                              (@                      @      2@                      @      @                      @      �?                      @                                      �?                              @                      �?      *@                      �?       @                               @                      �?                                      &@                       @                              @                                      1@                      �?     �\@                      �?      "@                              @                      �?      @                      �?      �?                      �?                                      �?                              @                             �Z@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJu�7hG        hNhG        hHKhIKhJh(h+K ��h-��R�(KK��hb�C               �?       @      @�t�bhVhghQC       ���R�hkKhlhoKh(h+K ��h-��R�(KK��hQ�C       �t�bK��R�}�(hKhyMhzh(h+K ��h-��R�(KM��h��B��         b                   �?T㥛���?�            �@       �                    "�@���n��?�           p�@       �                    -@�*���?=           �~@       5                    ��@��2'#r�?0           �}@                            #@��3L��?<             [@                          �H@��Wϊ�?              N@              	            Ɯ@�\ژW�?            �I@                           �?ףp=
�?             4@	       
                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �        
             1@                           @V��z4��?             ?@                           �?      �?              @                        `ff@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @                           @P���� �?             7@                           �?�a�a�?
             5@                           @���Q��?             @������������������������       �                     @������������������������       �                      @                           �?      �?             0@������������������������       �                     @                           �?B{	�%��?             "@                           t�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     "@!       2                   �2@VUUUU�?             H@"       /                    �?T�r
^N�?             E@#       .                   �E@�ͫ�gE�?             >@$       +                   �@@�8��8��?             8@%       (       	            ڢ@�ӭ�a��?	             2@&       '                     @      �?              @������������������������       �                     �?������������������������       �                     �?)       *       
             @      �?             0@������������������������       �                     �?������������������������       �                     .@,       -                    �?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @0       1       	            h�@r�q��?
             (@������������������������       �                      @������������������������       �                     $@3       4                   @F@r�q��?             @������������������������       �                     @������������������������       �                     �?6       Y                    �?ukL�v�?�            �v@7       @                    @y�����?1            @R@8       9       	            ��@��>��?            �E@������������������������       �                     <@:       ?       	            ��@���ĳ��?             .@;       <                    �?"pc�
�?	             &@������������������������       �                     �?=       >                    1@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?������������������������       �                     @A       L                    '@�������?             >@B       I                    �?�q�q�?	             (@C       H       
             -@և���X�?             @D       E                    �?z�G�z�?             @������������������������       �                     @F       G       	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @J       K                     @z�G�z�?             @������������������������       �                     �?������������������������       �                     @M       T       
             *@��Kh/�?             2@N       O                    �?��!pc�?             &@������������������������       �                     @P       S                    �?      �?             @Q       R       	            ;�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?U       X                    �?�$I�$I�?             @V       W                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @Z       �       	            h�@ �0����?�            0r@[       z                    �?M�Y�#�?p            �e@\       g                    �?��,�X�?=            �U@]       ^       	            H�@:ɨ��?            �@@������������������������       �                     5@_       f                    @r�q��?	             (@`       e                     @z�G�z�?             $@a       b                   �0@�����H�?             "@������������������������       �                     @c       d       
             +@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @h       i       	            p�@���_�?#            �J@������������������������       �                     1@j       m                    @���Kh�?             B@k       l       	            |�@      �?             @������������������������       �                     @������������������������       �                     �?n       o                 033�?     ��?             @@������������������������       �        
             2@p       s                    5@����S�?
             ,@q       r                    %@      �?              @������������������������       �                     �?������������������������       �                     �?t       u       	            V�@�8��8��?             (@������������������������       �                     @v       w                    $@z�G�z�?             @������������������������       �                     �?x       y                    @      �?             @������������������������       �                     �?������������������������       �                     @{       �                 ���@~�4_�g�?3             V@|       �                    �?�D����?0             U@}       �                    H�@�q�q�?            �C@~                           @��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@�       �       
            �3@      �?             8@�       �                    0@և���X�?             5@�       �                 ���@և���X�?
             ,@�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                 ���@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	            <�@��S���?            �F@�       �       	            4�@���7�?             6@������������������������       �                     4@�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     7@������������������������       �                     @�       �       
             -@+Jx��?S            @]@�       �                    5@ɢ4�N;�?<            @T@�       �       	            W�@l��
I��?             ;@�       �       
             %@P���Q�?
             4@������������������������       �                     .@�       �                    Ћ@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    �?����0�?,             K@�       �       	            �@      �?             4@������������������������       �                      @�       �       	            ��@r�q��?
             (@�       �       
             #@�q�q�?             @������������������������       �                     @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�       �       	            ��@�(��d��?             A@�       �       	            ��@؇���X�?             @�       �                    2�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    J@ 7���B�?             ;@������������������������       �                     7@�       �                    @      �?             @������������������������       �                     @������������������������       �                     �?�       �       
            �3@*O���?             B@�       �                    N@�;�;�?             :@�       �                 033�?`�Q��?             9@������������������������       �        	             *@�       �                    ,�@r�q��?	             (@�       �                    �?�8��8��?             @������������������������       �                      @�       �                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�       �                    �?ףp=
��?             $@������������������������       �                     @�       �                   �K@���Q��?             @������������������������       �                      @������������������������       �                     @�       �       
             @^Cy�5�?             3@�       �                   �1@      �?              @������������������������       �                     �?������������������������       �                     @�       �                    1@��!pc�?             &@�       �       	            ��@h/�����?             "@������������������������       �                      @�       �                    �?����X�?             @������������������������       �                     @�       �                    ^�@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�       E      	            ��@Z�L�$�?�            0r@�                          ��@���2��?w            �d@�                          '@�G�z��?;             T@�       �                    8@��ӭ�a�?3             R@�       �                 ���@ףp=
��?             >@�       �                    @�b��g�?             =@�       �                    ��@��Q��?	             $@������������������������       �                      @�       �                    @      �?              @�       �                    �?      �?             @������������������������       �                      @�       �                    %@      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @��uJ���?             3@�       �                    (@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    @     ��?             0@�       �       	            ��@�8��8��?             @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@������������������������       �                     �?�       �                 ����?.0�w¹�?             E@������������������������       �                     "@�       �                    �?8�#�(�?            �@@�       �       	            L�@tk~X��?             2@������������������������       �                     *@�       �                    �?���Q��?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       �       	            ��@VUUUUU�?
             .@������������������������       �                     @�                       033�?      �?             $@�                          $�@����X�?             @�                          �?r�q��?             @�       �                    �?�q�q�?             @������������������������       �                     �?                          "@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @                        �1@      �?              @      
                   0@0�����?             @      	                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?      :      
            �1@Ԁ�����?<            �U@                         �?�'}�'}�?3            �R@            	            �@VUUUUU�?	             .@������������������������       �                     @            	            `�@      �?             $@������������������������       �                     @������������������������       �                     @      )                   �?�������?*             N@                      ����?��S�r
�?             <@                      ����?�����H�?             "@            
             @r�q��?             @������������������������       �                     �?                         ʜ@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                         ��@��d����?             3@������������������������       �                     @      &                   �?6�h$��?             .@       %      	            ��@      �?              @!      "                   �@�q�q�?             @������������������������       �                     �?#      $      	            X�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @'      (                   Λ@؇���X�?             @������������������������       �                     �?������������������������       �                     @*      -                `ff�?      �?             @@+      ,                   r�@z�G�z�?             $@������������������������       �                      @������������������������       �                      @.      5                   �@��#��Z�?             6@/      4                pff�?�<ݚ�?             2@0      1                   �?      �?              @������������������������       �                     @2      3                   @z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@6      7                  �6@      �?             @������������������������       �                     �?8      9      	            ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @;      B                  �?@�q�q�?	             (@<      =      
            �2@�$I�$I�?             @������������������������       �                     @>      ?                033�?      �?             @������������������������       �                      @@      A                   �?      �?              @������������������������       �                     �?������������������������       �                     �?C      D      	            �@z�G�z�?             @������������������������       �                     @������������������������       �                     �?F      G                   @8��d�?I             _@������������������������       �                      @H      ]                  �B@�t`�4 �?H            �^@I      X      
            �2@h�˹�?,             S@J      M                   �?@�j;��?(            �Q@K      L                  �3@�(\����?             D@������������������������       �                    �C@������������������������       �                     �?N      S                   ��@�חF�P�?             ?@O      R                  �>@���Q��?             $@P      Q                   ��@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @T      W                   �?���N8�?             5@U      V      	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        
             3@Y      Z                   @���Q��?             @������������������������       �                     �?[      \                   �?      �?             @������������������������       �                     �?������������������������       �                     @^      a                   4�@�nkK�?             G@_      `                   ��@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                    �B@c      �                   -@*"�+��?           ��@d      �                   �?�(�4g��?y           ��@e      �                   @��� Ce�?<            �V@f      s                   %@L�t��>�?$             K@g      j                   �?��ˠ�?             &@h      i      	            I�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @k      p                   �?VUUUUU�?             @l      m                   @      �?             @������������������������       �                      @n      o                   !@      �?              @������������������������       �                     �?������������������������       �                     �?q      r                   �?      �?              @������������������������       �                     �?������������������������       �                     �?t      �                   �?ZJj�?            �E@u      |                   �?(������?             3@v      w                  �K@ףp=
�?             $@������������������������       �                     @x      y                   @z�G�z�?             @������������������������       �                     @z      {                  @M@      �?              @������������������������       �                     �?������������������������       �                     �?}      ~      
             @x�5?,�?             "@������������������������       �                      @      �      	            �@0�����?             @������������������������       �                     @�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �@9��8���?             8@�      �      	            v�@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�      �      
             3@�(ݾ�z�?             *@�      �                   �@VUUUUU�?             "@�      �      
             /@z�G�z�?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �@      �?             @������������������������       �                      @�      �                @33�?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @�      �                   @\��"e��?             B@�      �                   D�@#AM�h��?             :@�      �      
             &@$I�$I��?             ,@�      �                   /@X�<ݚ�?             "@������������������������       �                      @�      �                   ��@����X�?             @�      �                  �3@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                hff�?�Q����?             @������������������������       �                     �?�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @�      �                  �@@9��8���?	             (@�      �                  �5@z�G�z�?             @������������������������       �                     @�      �                ����?      �?              @������������������������       �                     �?������������������������       �                     �?�      �      	            
�@և���X�?             @������������������������       �                     @������������������������       �                     @�      �                   9@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@�      �                   @]��z��?=           �@�      �      	            ϣ@���Q��?             D@�      �                   @{�G�z�?
             4@�      �      	            ��@      �?              @������������������������       �                     @�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @�      �                   @�q�q�?             (@�      �                  @F@������?             @�      �                   @      �?             @������������������������       �                     �?�      �                  �7@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @�      �      
             @P���Q�?
             4@�      �                  @@@      �?              @������������������������       �                     @�      �                   ��@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�      -      	            ܡ@B�7����?)           }@�      �      	            |�@�'n�N�?�            @p@�      �                   �?���}<S�?M            �\@�      �      	            `�@      �?             @������������������������       �                      @������������������������       �                      @�      �                   @���l��?I            �[@�      �      	            0�@���!pc�?             &@�      �                   �?�����H�?             "@�      �                  �E@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                  �O@P���Q�?A             Y@�      �                   >@`�(c�??            �X@������������������������       �        #            �K@�      �                ����?Du9iH��?            �E@�      �                033�?�LQ�1	�?             7@�      �      
            �2@�X�<ݺ?
             2@������������������������       �        	             1@������������������������       �                     �?�      �                   @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     4@������������������������       �                      @�                         @T�ǹ�#�?]             b@�      �                ����?V�h3��?O            @^@�      �                   �?��y�):�?             9@�      �      	            >�@
ц�s�?
             *@�      �      
             /@���Q��?             $@�      �      	            ��@      �?              @������������������������       �                      @������������������������       �                     @������������������������       �                      @������������������������       �                     @�      �      
             +@�q�q�?             (@�      �                   �?      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                     @�                         �?�����*�?@             X@�      
                   @0E�f���?            �G@�      	                   &�@�n_Y�K�?            �C@�      �                   ��@��Coul�?            �B@������������������������       �                      @�      �                   @"	��p�?             =@������������������������       �                      @�                         +@�5��?             ;@�      �                   @`�Q��?             9@�      �                   �?      �?              @������������������������       �                     @������������������������       �                     @                         @K@�"�O�|�?             1@            	            ��@      �?
             0@                         @      �?              @������������������������       �                     �?            	            ԕ@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @            	            D�@�2�|�&�?#            �H@                         @��
ц��?
             *@                         @���Q��?             $@������������������������       �                     @                      ���@؇���X�?             @������������������������       �                     @                         l�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                         @�8��8��?             B@������������������������       �        	             0@                      pff�?R���Q�?             4@������������������������       �                     "@                         @���!pc�?
             &@������������������������       �                     @������������������������       �                      @                      ����?9��8���?             8@������������������������       �                     @      "                   3@���(\��?             4@       !                   �?؇���X�?             @������������������������       �                     �?������������������������       �                     @#      *      
             1@8�Z$���?
             *@$      %                pff@B{	�%��?             "@������������������������       �                     @&      '                   �?VUUUUU�?             @������������������������       �                     �?(      )                   %@      �?              @������������������������       �                     �?������������������������       �                     �?+      ,                  �9@      �?             @������������������������       �                     �?������������������������       �                     @.      /                   @�/Sh�'�?            �i@������������������������       �                     (@0      S                   Đ@pɂ��?z             h@1      N                   @6?,R��?1             R@2      =                   �?L�.�o�?$            �I@3      6                ����?      �?             8@4      5      	            ��@      �?              @������������������������       �                     @������������������������       �                     @7      :                   @     ��?             0@8      9      	            ��@      �?              @������������������������       �                     @������������������������       �                     @;      <                   �?      �?              @������������������������       �                      @������������������������       �                     @>      M                   @F&K:�m�?             ;@?      L                   @p=
ףp�?             4@@      G                   �@���Q��?             .@A      B                   �?�Q����?             @������������������������       �                     �?C      D                   @      �?             @������������������������       �                      @E      F                   N@      �?              @������������������������       �                     �?������������������������       �                     �?H      I                   \�@ףp=
�?             $@������������������������       �                     @J      K                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @O      P      
            �0@؇���X�?             5@������������������������       �                     (@Q      R                   �?�q�q�?             "@������������������������       �                     @������������������������       �                     @T      {      
            �1@��,?S�?I            @^@U      `                   ș@���c��?=            �W@V      _      	            �@Riv����?$             M@W      Z                   �?X�Cc�?             ,@X      Y                   l�@���Q��?             @������������������������       �                     @������������������������       �                      @[      \                033�?�q�q�?             "@������������������������       �                      @]      ^                   @؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     F@a      d                   @��+��?            �B@b      c                ����?r�q��?             @������������������������       �                     @������������������������       �                     �?e      r                    @`՟�G��?             ?@f      k      
             "@�X����?             6@g      j                   �@r�q��?             @h      i                ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @l      q                   ��@      �?
             0@m      p      	            �@��S�ۿ?	             .@n      o      
             /@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?s      z                   �?�<ݚ�?             "@t      y                   �?����X�?             @u      x                   �?r�q��?             @v      w                   @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?������������������������       �                      @|      }                   +@ ��WV�?             :@������������������������       �        
             6@~                         �?      �?             @������������������������       �                     �?������������������������       �                     @�      �                   �?�R�h���?�            �k@�      �      	            Ȥ@      �?             0@�      �                   D�@      �?              @������������������������       �                     @�      �                  �0@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @�      �                  �0@h�V�w<�?~            �i@�      �                   @kN¾��?$            �L@�      �      	            Ȟ@&�9�٫�?            �B@�      �                   �?�<ݚ�?             "@������������������������       �                     @�      �      
             .@      �?             @������������������������       �                      @������������������������       �                      @�      �                   @ܶm۶m�?             <@�      �      	            A�@��ͦ-��?             ;@�      �                   �? �q�q�?             8@������������������������       �                     *@�      �                   @�C��2(�?             &@������������������������       �                     "@�      �      	            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   ��@��Q���?             4@�      �                   ��@P�|�@�?             1@�      �                   @      �?              @������������������������       �                      @�      �      
             !@      �?             @������������������������       �                     @�      �                033�?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  �C@�n���?             "@�      �                   1@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                     @�      �                   @4��!j�?Z            �b@�      �                   ��@��FZ���?;            @X@�      �                   �?������?%             L@�      �      	            �@�mM`���?             7@������������������������       �        
             *@�      �      	            k�@p=
ףp�?	             $@������������������������       �                     @�      �                   K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   0�@6YE�t�?            �@@�      �      
             +@b���i��?             &@�      �                033@������?             @�      �                   �?�Q����?             @�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �      
             @�eP*L��?             6@�      �                   3@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   2@�G�z��?
             4@������������������������       �                     �?�      �      	            ,�@�}�+r��?	             3@������������������������       �                     �?������������������������       �                     2@�      �                   '@��t���?            �D@�      �                   �?L�6�#��?             ?@�      �                  �1@{�G�z�?             .@�      �      	            N�@:/����?             @�      �                  �F@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                      @�      �      	            *�@     ��?
             0@�      �                   @8�Z$���?             *@�      �                   �?�8��8��?             (@�      �                  @A@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     �?�      �                   K@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   @ףp=
�?             $@�      �                   .@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                   �?��b�,��?            �J@�      �      	            ��@VUUUUU�?             8@�      �      	            H�@�r����?             .@�      �      	            �@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @�      �                   @�n���?             "@�      �                  �A@�Q����?             @�      �      	            |�@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �                   �?      �?             @�      �                @33�?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�      �      
             "@ܷ��?��?             =@�      �                `ff @��8��8�?             (@�      �                   �@�z�G��?             $@�      �                   ,�@      �?              @������������������������       �                     @�      �                   2@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                      @�                          �?�������?	             1@�      �                   �?؇���X�?             @������������������������       �                     @������������������������       �                     �?                         �?H�z�G�?             $@                         ؝@r�q��?             @������������������������       �                     @������������������������       �                     �?                          @      �?             @������������������������       �                     @������������������������       �                     �?�t�b�X-     h�h(h+K ��h-��R�(KMKK��hb�B�`       0z@     �y@     �w@     �x@      h@     `i@     �h@     �g@     �a@     �a@     �`@     �R@     �a@      a@      `@     @P@      9@      =@      G@       @      2@      4@      2@      @      2@      &@      2@      @      2@       @                      �?       @                      �?                                       @                      1@                                      "@      2@      @              @       @                      @       @                      @                                       @                      @                              @      0@      @              �?      0@      @                       @      @                              @                       @                      �?      ,@      �?                      @                      �?      @      �?              �?              �?              �?                                              �?                      @                       @                              "@                      @      "@      <@      @      @      @      ;@      @      @       @      1@      @      �?       @      1@      @      �?       @      .@              �?      �?                      �?                                      �?                              �?      .@                      �?                                      .@                               @      @                       @                                      @      @                                       @      $@                       @                                      $@                      @      �?                      @                                      �?             �]@     �Z@     �T@     �L@      B@      (@      4@      @      <@       @      "@      @      <@                                       @      "@      @               @      "@                      �?                              �?      "@                              "@                      �?                                              @       @      $@      &@      �?      @       @              �?      @      @                      �?      @                              @                      �?      �?                      �?                                      �?                       @                                      @              �?                              �?              @                      @       @      &@              �?      �?      "@                              @              �?      �?       @                      �?       @                      �?                                       @              �?                              @      �?       @              @      �?                              �?                      @                                               @             �T@     �W@      O@      J@     �T@     �V@      �?              F@     �D@      �?              7@      $@                      5@                               @      $@                       @       @                      �?       @                              @                      �?       @                      �?                                       @                      �?                                       @                      5@      ?@      �?              1@                              @      ?@      �?              @      �?                      @                                      �?                      �?      >@      �?                      2@                      �?      (@      �?              �?      �?                              �?                      �?                                      &@      �?                      @                              @      �?                      �?                              @      �?                              �?                      @                      C@      I@                      A@      I@                      *@      :@                      �?      ,@                      �?                                      ,@                      (@      (@                      (@      "@                      @       @                      �?      @                      �?                                      @                      @      �?                      @                                      �?                      @      �?                      @                                      �?                              @                      5@      8@                      5@      �?                      4@                              �?      �?                              �?                      �?                                      7@                      @                                      @     �N@      J@              �?      B@      F@                      3@       @                      3@      �?                      .@                              @      �?                      @                                      �?                              @              �?      1@      B@                      $@      $@                       @                               @      $@                       @      @                              @                       @      �?                       @                                      �?                              @              �?      @      :@              �?      @                      �?      �?                              �?                      �?                                      @                              �?      :@                              7@                      �?      @                              @                      �?                      @      9@       @              �?      6@      @              �?      6@       @                      *@                      �?      "@       @              �?      @       @                               @              �?      @                      �?                                      @                              @                                      �?               @      @      @                              @               @      @                       @                                      @                      @      @      "@                      �?      @                      �?                                      @              @      @       @               @      @       @               @                                      @       @                      @                               @       @                       @                                       @               @                     �H@     �O@      P@     �\@     �H@     �O@     �I@      @      B@      3@      8@      �?      A@      ,@      7@      �?      @      @      0@      �?      @      @      0@      �?      @      @      @               @                              �?      @      @                      @      @                               @                      @      �?                              �?                      @                      �?      �?                      �?                                      �?                      @      �?      *@      �?       @      �?                              �?                       @                               @              *@      �?       @              @      �?       @                      �?       @                                                      �?                      @                              $@                      �?                      ;@       @      @              "@                              2@       @      @              *@      @       @              *@                                      @       @                      @      �?                              �?                      @                                      �?              @      @      @              @                                      @      @                      @       @                      @      �?                       @      �?                      �?                              �?      �?                      �?                                      �?                      @                                      �?                              @               @      @      �?              �?      @      �?              �?              �?                              �?              �?                                      @                      �?                              *@      F@      ;@      @      "@      E@      7@      �?      @      @      @              @                                      @      @                      @                                      @              @     �B@      2@      �?      �?      ,@      (@      �?               @      �?                      @      �?                      �?                              @      �?                              �?                      @                              @                      �?      @      &@      �?              @                      �?       @      &@      �?      �?       @      @              �?       @                              �?                      �?      �?                      �?                                      �?                                      @                              @      �?                              �?                      @              @      7@      @               @       @                       @                                       @                      �?      .@      @                      ,@      @                      @      @                              @                      @      �?                      @                                      �?                      $@                      �?      �?       @              �?                                      �?       @                      �?                                       @              @       @      @       @               @      @      �?                      @                       @      �?      �?               @                                      �?      �?                              �?                      �?              @                      �?      @                                                      �?                      *@     �[@                       @                              &@     �[@                      "@     �P@                      @     @P@                      �?     �C@                             �C@                      �?                              @      :@                      @      @                      @       @                               @                      @                                      @                      �?      4@                      �?      �?                      �?                                      �?                              3@                      @       @                              �?                      @      �?                              �?                      @                               @      F@                       @      @                              @                       @                                     �B@     `l@     �i@     @f@      j@     �e@      a@     @\@     �e@     �@@      2@      5@      2@      :@      (@      @      (@      �?      @      �?      @              �?              @              �?                                              @      �?      @      �?      �?              @              �?               @                              �?              �?                              �?              �?                      �?              �?                              �?              �?                              9@       @      @      @      ,@       @              @      "@      �?                      @                              @      �?                      @                              �?      �?                              �?                      �?                              @      �?              @                               @      @      �?              �?      @                                      �?              �?              �?                                              �?      &@      @      @      @      "@       @                      "@                                       @                       @      @      @      @      �?      �?      @      @                      �?      @                      �?      �?                      �?                                      �?                              @      �?      �?       @                               @              �?      �?                      �?                                      �?                      �?      @                      �?                                      @                      @      @      1@      @      @      @       @      @      @      @      @                      @      @                               @                      @       @                      �?       @                      �?                                       @                      @                      @      �?      �?                              �?              @      �?                              �?                      @                              @              @      @      @                      �?      @                              �?                      �?      �?                                                      �?                      @      @                      @                                      @                      "@      �?                              �?                      "@             `a@     �]@      W@     �c@       @       @      @      3@       @       @      @                      @      �?                      @                              @      �?                              �?                      @                       @      �?      @              @      �?      @              @      �?                      �?                               @      �?                              �?                       @                                              @              @                                              �?      3@                      �?      @                              @                      �?      @                      �?                                      @                              (@     ``@     �[@     �U@      a@     ``@     �Z@      7@             @Z@      $@                       @       @                       @                                       @                     �Y@       @                       @      @                       @      �?                      @      �?                      @                                      �?                      @                                       @                     �W@      @                     �W@      @                     �K@                              D@      @                      4@      @                      1@      �?                      1@                                      �?                      @       @                      @                                       @                      4@                                       @                      :@      X@      7@              0@      V@      1@               @      ,@      @              @      @      @              @      @                       @      @                       @                                      @                       @                                              @              @       @                      @      @                      @                                      @                              @                       @     �R@      ,@               @      A@      &@               @      :@      &@               @      :@      "@                       @                       @      2@      "@                               @               @      2@      @               @      2@      @                      @      @                              @                      @                       @      ,@      �?               @      ,@                       @      @                      �?                              �?      @                              @                      �?                                       @                                      �?                               @                               @                       @                      @      D@      @              @      @                      @      @                              @                      @      �?                      @                              �?      �?                      �?                                      �?                              @                             �@@      @                      0@                              1@      @                      "@                               @      @                              @                       @                      $@       @      @                              @              $@       @       @              @              �?                              �?              @                              @       @      �?              �?      @      �?                      @                      �?      �?      �?                              �?              �?      �?                      �?                                      �?                      @      �?                              �?                      @                                      @      P@      a@                              (@              @      P@     @_@              @     �A@     �@@              @      @@      .@              @      .@      @                      @      @                      @                                      @              @      &@       @              @      @                      @                                      @                              @       @                               @                      @                      �?      1@      "@              �?      $@      "@              �?      $@      @              �?      �?      @                      �?                      �?              @                               @              �?              �?              �?                                              �?                      "@      �?                      @                               @      �?                       @                                      �?                              @                      @                              @      2@                              (@                      @      @                              @                      @                              =@      W@                      <@     �P@                      "@     �H@                      "@      @                      @       @                      @                                       @                      @      @                               @                      @      �?                      @                                      �?                              F@                      3@      2@                      @      �?                      @                                      �?                      ,@      1@                      @      .@                      @      �?                      �?      �?                      �?                                      �?                      @                               @      ,@                      �?      ,@                      �?      @                              @                      �?                                      &@                      �?                              @       @                      @       @                      @      �?                       @      �?                              �?                       @                              @                                      �?                       @                              �?      9@                              6@                      �?      @                      �?                                      @     �K@     @Q@     @P@      A@      @       @       @       @      @       @       @              @                                       @       @                               @                       @                                               @     �I@     �P@     �O@      :@       @      ,@      :@      "@       @       @      7@      @       @      @                              @                       @       @                               @                       @                                      �?      7@      @              �?      7@      @              �?      7@                              *@                      �?      $@                              "@                      �?      �?                      �?                                      �?                                      @                              �?      @      @      @      @      @      @      @      @      @      @              �?               @                      @      �?              �?      @                                      �?              �?              �?                                              �?       @              @      @       @              @                              @               @                                                      @              @                     �E@     �J@     �B@      1@      6@     �E@      8@       @      2@      =@      @      @      *@      @      �?       @      *@                                      @      �?       @              @                                      �?       @                               @                      �?              @      6@      @       @      @      @      @      �?              @      @      �?              @      �?      �?              @              �?              @                                              �?                      �?                               @              @                              �?      3@      �?      �?              �?      �?                              �?                      �?                      �?      2@              �?                              �?      �?      2@                      �?                                      2@                      @      ,@      3@      @      @      *@      $@      @       @       @       @      @       @       @              @       @       @                       @                                       @                                              @                       @               @      &@       @      �?       @      &@                      �?      &@                      �?      @                      �?                                      @                              @                      �?                                               @      �?                       @                                      �?              �?      "@                      �?      @                              @                      �?                                      @              5@      $@      *@      "@      *@      @      @      @      *@       @                      @       @                      @                                       @                       @                                       @      @      @              �?      @      �?              �?      @                      �?                                      @                                      �?              �?      �?       @              �?               @                               @              �?                                      �?               @      @      "@      @       @      @      @                      @      @                      �?      @                              @                      �?       @                      �?                                       @                       @                       @                              @      @       @      @      @              �?              @                                              �?                      @      �?      @                      �?      @                              @                      �?                      @              �?              @                                              �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ��!XhG        hNhG        hHKhIKhJh(h+K ��h-��R�(KK��hb�C               �?       @      @�t�bhVhghQC       ���R�hkKhlhoKh(h+K ��h-��R�(KK��hQ�C       �t�bK��R�}�(hKhyM�hzh(h+K ��h-��R�(KM���h��B8�         �                    �?u���?�            �@       �                   �F@D�d��?�            �x@       &                    @�8�����?�            �q@              	            ��@�|/D �?#             M@                           .@�w�AV�?            �E@                           &@Y�����?             &@       
                    @      �?             @       	                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @              	            ��@      �?             @@������������������������       �                     @                          �C@��)x9�?             <@                           �?P���� �?             7@                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           @P���Q�?	             4@������������������������       �                     (@                            @      �?              @                           @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                           �?{�G�z�?             @                           @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @        %                    @z�G�z�?
             .@!       $                   �4@$�q-�?	             *@"       #                    �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     "@������������������������       �                      @'       �                    !@��X��?�             l@(       =                    %@���h��?{            �g@)       4                    @j����?             =@*       /                    �?���k���?             &@+       .                 ���@����X�?             @,       -       
             "@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?0       1                     @      �?             @������������������������       �                     �?2       3       	            l�@�q�q�?             @������������������������       �                      @������������������������       �                     �?5       6       	            �@���[���?             2@������������������������       �                     @7       8                    �?�θ�?
             *@������������������������       �                     @9       :                    �?և���X�?             @������������������������       �                      @;       <                    $�@���Q��?             @������������������������       �                      @������������������������       �                     @>       K                    +@{�G��?f             d@?       @                 033�?�˹�m��?             3@������������������������       �                     @A       J                 ����?     ��?	             0@B       G                    '@�<ݚ�?             "@C       F                    %@{�G�z�?             @D       E                    ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @H       I                    )@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @L       g       
             )@��R�/z�?[            �a@M       ^                    x�@'&��|��?,            �P@N       S       	            ��@�u�Ë��?#             K@O       R                    @���7�?             6@P       Q       	            ^�@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     0@T       U                    �?     P�?             @@������������������������       �                      @V       ]       	            ��@�q�q�?             8@W       \                    @��(\���?	             $@X       Y                    @�����H�?             "@������������������������       �                     @Z       [       	            {�@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     ,@_       `                    ��@��WV��?	             *@������������������������       �                     @a       d                    �?�$I�$I�?             @b       c                    ڞ@z�G�z�?             @������������������������       �                     �?������������������������       �                     @e       f                    �@      �?              @������������������������       �                     �?������������������������       �                     �?h       �                    @qD���?/            �R@i       v       	            ��@4�����?(             O@j       q                 `ff�?��X��?             <@k       n                     @;�;��?             *@l       m                    @r�q��?             @������������������������       �                     �?������������������������       �                     @o       p                   �6@����X�?             @������������������������       �                      @������������������������       �                     @r       s                    @H�7�&��?             .@������������������������       �                     �?t       u       	            6�@؇���X�?             ,@������������������������       �                      @������������������������       �        
             (@w       z                 033�?��.k���?             A@x       y                   �A@؇���X�?             @������������������������       �                     @������������������������       �                     �?{       |       	            k�@��}*_��?             ;@������������������������       �                     @}       ~                    ��@�GN�z�?             6@������������������������       �                     @       �                    0�@�KM�]�?             3@�       �                 ���@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     *@�       �       	            7�@�8��8��?             (@������������������������       �                     $@�       �                    '@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?���Ze��?            �A@�       �       
             &@�n���?	             2@������������������������       �                     @�       �                    -@�؉�؉�?             *@������������������������       �                      @�       �                    �@�Q����?             @�       �                    �?      �?             @�       �                    $@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�       �                    @|�/��>�?
             1@������������������������       �                      @�       �                    /@��E���?             "@�       �       	            ̎@0�����?             @������������������������       �                     �?�       �                    A@r�q��?             @������������������������       �                     @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?�       �       
            �3@#��
��?C            �[@�       �                    �?�O��n�?;             Y@�       �                    �?�KL���?            �B@������������������������       �                      @�       �                    ��@��@z��?            �A@�       �                    �?E3����?             ;@�       �       
             @     ��?
             0@������������������������       �                     @�       �                    J@p=
ףp�?             $@�       �                    ��@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     @�       �                 ����?"pc�
�?             &@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�       �                    �?      �?              @�       �                    �?      �?             @������������������������       �                      @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �       
              @&)��a�?%            �O@�       �                    �?     ��?             0@�       �       	            @�@      �?              @������������������������       �                     @������������������������       �                     @�       �       	            /�@      �?              @�       �                    �?�q�q�?             @������������������������       �                     �?�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    �?��9���?            �G@�       �                   �L@�lO���?
             3@�       �       	            �@;�;��?             *@������������������������       �                     @�       �                    X�@����X�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�       �       	            ��@x9/���?             <@�       �       
             /@�lO���?
             3@�       �                    @8�Z$���?             *@�       �                   �K@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                   �H@�����H�?             "@������������������������       �                     �?������������������������       �                      @�       �                    !@���(\��?             $@�       �                    �?      �?              @�       �                     @VUUUUU�?             @������������������������       �                     �?�       �       	            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�       �                    ��@      �?              @������������������������       �                     �?������������������������       �                     �?�       ^                   �?��]`���?�           ��@�       �                   ��@_3UYp��?�           8�@�       �                   >�@z%�V�(�?�            pv@�                          @��|�`a�?�             u@�             
             /@��j�e{�?:            �Z@�       �       
             @��&�v�?/            �V@�       �                    @�X�C�?             ,@�       �                    5@���k���?             &@������������������������       �                      @�       �                 033�?�<ݚ�?             "@������������������������       �                      @������������������������       �                     @������������������������       �                     @�                       hff @;�lO�?)             S@�       �       	            ��@�F�P�?!             O@������������������������       �        	             0@�       �                 ����?ԛ���7�?             G@�       �                    �?��8��8�?             (@������������������������       �                      @�       �                    F@H�z�G�?             $@�       �                    (@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�                          ��@�������?             A@�                          @�h��U�?            �@@�                          !@��eP*L�?             6@                       pff�?��S�ۿ?             .@                         �?r�q��?             @                         @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     "@            	            �@:/����?             @������������������������       �                     @	      
                   �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     &@������������������������       �                     �?                         @������?             ,@                         @z�G�z�?             @������������������������       �                      @                         ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         ��@�n���?             "@������������������������       �                     @                         �?���Q��?             @������������������������       �                     �?                         �@      �?             @������������������������       �                     �?������������������������       �                     @            	            ��@     ��?             0@������������������������       �                     *@                         @�q�q�?             @������������������������       �                     �?������������������������       �                      @       �      
            �3@ �v)�?�?�            �l@!      ~                   @d}h�-�?�             l@"      ?                   �@ \��M�?T             a@#      &      
             @(�כbv�?!            �J@$      %      	            M�@؇���X�?             @������������������������       �                     �?������������������������       �                     @'      (      	            ��@���?             G@������������������������       �                     *@)      .                  �7@'�`de�?            �@@*      +                   @ףp=
�?             $@������������������������       �                     @,      -      	            ��@      �?             @������������������������       �                     �?������������������������       �                     @/      2                   X�@h�d0ܩ�?             7@0      1                   4�@؇���X�?             @������������������������       �                     �?������������������������       �                     @3      :                   �?     ��?
             0@4      9                   �?r�q��?             @5      8                   �?z�G�z�?             @6      7      	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     �?;      >                  @I@H�z�G�?             $@<      =                  �8@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @@      w                   @�Q�@��?3            �T@A      P                   @     ��?)             P@B      E      
             @2�tk~X�?             2@C      D                   &@      �?             @������������������������       �                     @������������������������       �                     �?F      K                   @������?
             ,@G      H      	            �@      �?              @������������������������       �                     @I      J                   �?      �?              @������������������������       �                     �?������������������������       �                     �?L      O                   !@�q�q�?             @M      N                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?Q      V                   ��@
,UP���?             G@R      S                   C@�8��8��?             (@������������������������       �                     "@T      U      	            �@�q�q�?             @������������������������       �                     �?������������������������       �                      @W      f                   �?�7�
t��?             A@X      Y      
             @N��)x9�?
             ,@������������������������       �                     @Z      _                   �?�x?r���?             &@[      ^                   @{�G�z�?             @\      ]      	            �@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @`      a      
             /@VUUUUU�?             @������������������������       �                     @b      c                   ��@VUUUUU�?             @������������������������       �                     �?d      e                   @      �?              @������������������������       �                     �?������������������������       �                     �?g      n      
              @�Q����?             4@h      k                   ��@p=
ףp�?             $@i      j                   �?���Q��?             @������������������������       �                      @������������������������       �                     @l      m                   8@z�G�z�?             @������������������������       �                     �?������������������������       �                     @o      v                   ��@p=
ףp�?             $@p      u                   @B{	�%��?             "@q      r                   �?      �?              @������������������������       �                     @s      t                   "@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     �?x      {                   �?ԍx�V�?
             3@y      z                   F@�t����?             1@������������������������       �                     .@������������������������       �                      @|      }                   f�@      �?              @������������������������       �                     �?������������������������       �                     �?      �                   @�9����?>             V@�      �      	            ��@"pc�
�?            �@@�      �      
             @����X�?             @�      �                   �@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�      �                   +@ ��WV�?             :@�      �                   )@�C��2(�?             &@������������������������       �                     "@�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     .@�      �      
            �1@�"�����?*            �K@�      �      	            .�@VUUUU��?&             H@������������������������       �                     .@�      �                  �0@�x?r���?            �@@�      �                  �I@�p=
ף�?             4@�      �      
             +@      �?             0@�      �                   �?j�V���?	             &@�      �                   �?{�G�z�?             @�      �      
             $@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   ܊@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �?{�G�z�?             @������������������������       �                      @�      �                   2�@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?�      �                   .@�	j*D�?
             *@������������������������       �                     @�      �                   :�@���Q��?             $@�      �                  �1@z�G�z�?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                ��� @؇���X�?             @������������������������       �                     �?������������������������       �                     @�      �                   .@      �?             @������������������������       �                      @�      �                   �?      �?             @������������������������       �                      @�      �      	            @      �?              @������������������������       �                     �?������������������������       �                     �?�      �      	            �@8����?             7@������������������������       �                     0@������������������������       �                     @�                        �@@    ���?�             p@�      �                    �@��g�L��?\            �`@�      �                   ��@�z�G!�?2             T@�      �                   )@j�6�i�?'             N@�      �                ����?_�_��?            �A@�      �                   �?0�����?             @�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �      	            b�@      �?             <@�      �                   �?�t����?	             1@������������������������       �                     @�      �      	            ��@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�      �                   @��!pc�?             &@�      �                ����?0�����?             @������������������������       �                     �?�      �                pff@r�q��?             @������������������������       �                     @�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @�      �                ���@^K�=��?             9@�      �                ����?�}2��?             1@�      �                   �?pƵHP�?
             *@�      �                   �?z�G�z�?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                   �?      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �                   @      �?              @�      �                   @      �?             @�      �      
             @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   �?>
ףp=�?             4@�      �                   �@
ףp=
�?             @�      �                    @VUUUUU�?             @������������������������       �                     �?�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                   @��S�ۿ?             .@������������������������       �                     �?������������������������       �                     ,@�             	            �@^�vD'0�?*            �K@�      �                ���@r�q��?             8@�      �                   @     ��?             0@�      �                   ��@@4և���?             ,@�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �        	             (@������������������������       �                      @�      �                   �?      �?              @������������������������       �                     �?�      �                   0@؇���X�?             @������������������������       �                     @������������������������       �                     �?      
                   N�@���@M^�?             ?@      	      	            2�@R�}e�.�?             :@                         *@P���Q�?             4@                         &@ףp=
�?             $@������������������������       �                      @                         ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@������������������������       �                     @������������������������       �                     @                         ��@��/��n�?T            @^@            
             @D>�Q�?             :@������������������������       �                     "@                         �?��\���?             1@                         ��@X�<ݚ�?             "@            
             @�q�q�?             @������������������������       �                      @                      ����?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @                      `ff�?      �?              @            
             *@      �?              @������������������������       �                     �?������������������������       �                     �?                         �?r�q��?             @                        @I@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @       9                   @�՘���?D            �W@!      .      	            �@�d��)�?             �F@"      )                   @w���<�?             ?@#      (                   �?~h����?	             ,@$      '      	            L�@��8��8�?             (@%      &      	            @r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @*      +                   �?8߄*�u�?             1@������������������������       �                     �?,      -      	            `|@      �?
             0@������������������������       �                     �?������������������������       �        	             .@/      2                   @և���X�?             ,@0      1                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @3      4                   �?�<ݚ�?             "@������������������������       �                     �?5      6      
             +@      �?              @������������������������       �                     @7      8                ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @:      ?      
             @�.n���?$             I@;      <                   @      �?             @������������������������       �                     @=      >                   @      �?              @������������������������       �                     �?������������������������       �                     �?@      O                  @G@      �?             F@A      D                   �?8��8���?             8@B      C      
             +@�q�q�?             @������������������������       �                      @������������������������       �                     �?E      L                   @�&%�ݒ�?             5@F      K      	            ��@�eP*L��?             &@G      J      	            ��@r�q��?             @H      I                  �D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @M      N                ���@ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?P      ]                   @�G�z��?             4@Q      X                  �L@0��b�/�?             .@R      S      	            ��@��ˠ�?	             &@������������������������       �                     @T      U      	            ��@0�����?             @������������������������       �                     �?V      W                   @r�q��?             @������������������������       �                     �?������������������������       �                     @Y      \      
             !@      �?             @Z      [                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @_      h                   ��@�bն��?m           ��@`      g                033@���,�?             C@a      b      	            ܜ@��\���?             A@������������������������       �                     =@c      f                   �?�Q����?             @d      e                   �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @i                         �?rLB�W��?\           X�@j      �                   @Rn�?���?�            pr@k      �                   @x�����?x            �g@l      {                   �?$I�$I��?G             \@m      t                  �@@�p9W���?             3@n      o                   @z�G�z�?             $@������������������������       �                     @p      s                033�?�q�q�?             @q      r                  �0@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @u      x                   �?x�5?,�?             "@v      w                   �@z�G�z�?             @������������������������       �                     �?������������������������       �                     @y      z                   #@      �?             @������������������������       �                     @������������������������       �                     �?|      �                    @����C��?;            @W@}      �                   @�q�q�?             "@~                         �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �      	            ��@ܶm۶m�?5             U@�      �      
             #@�P�*�?             ?@�      �                   (@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?�      �      
             +@�q�q�?             2@������������������������       �                     @�      �                  �B@��
ц��?	             *@�      �                   �?؇���X�?             @�      �      	            ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �      
             #@�+����?#            �J@�      �                   ��@ �o_��?             9@�      �      	            b�@؇���X�?             5@������������������������       �                     @������������������������       �                     2@������������������������       �                     @�      �                   @�r
^N��?             <@�      �                   0�@>F?�!��?             5@������������������������       �                      @�      �      
             /@�S����?
             3@�      �      	            �@�z�G��?             $@������������������������       �                     @������������������������       �                     @������������������������       �                     "@������������������������       �                     @�      �                   �?��ײ���?1            �S@�      �                   @�m۶m��?             <@�      �      
             !@���Q��?             .@������������������������       �                     @�      �                   ��@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�      �      
             &@�؉�؉�?             *@������������������������       �                     "@�      �      	             �@      �?             @������������������������       �                     �?������������������������       �                     @�      �      	            ��@��Z�-�?"            �I@�      �                   6@     @�?             @@�      �                   �?      �?             (@������������������������       �                     "@������������������������       �                     @�      �                   �@
ףp=
�?             4@�      �      	            ��@�n_Y�K�?             *@������������������������       �                     @������������������������       �                      @�      �                ����?և���X�?             @������������������������       �                     @������������������������       �                     @�      �      	            �@�KM�]�?             3@�      �                  �L@���Q��?             @�      �                   �?�q�q�?             @������������������������       �                     �?�      �      	            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     ,@�      �                   �?/y0��k�?=             Z@�      �      	            ��@L�t��>�?             ;@�      �                   (@H�z�G�?             4@�      �                   x�@     ��?	             0@�      �                   @      �?              @������������������������       �                     @�      �                   �?      �?             @�      �                   !@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @�      �      
             3@      �?             @������������������������       �                     @������������������������       �                     �?�      �                  �H@؇���X�?             @������������������������       �                     @������������������������       �                     �?�      �                   @D�+ṗ�?-            @S@�      �                   �?9��8���?             8@�      �      	            !�@"pc�
�?             &@������������������������       �                     @�      �      
             @      �?              @������������������������       �                     �?�      �                   (@؇���X�?             @������������������������       �                     �?������������������������       �                     @�      �                   �?pƵHP�?             *@�      �                ����?      �?              @������������������������       �                     @�      �      	            ޝ@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @�      	                033@�2s��?            �J@�      �                   @W�+���?            �G@������������������������       �                     @�      �                   #@�G�z�?             D@�      �                ���@)O���?             2@�      �      
             #@     @�?
             0@�      �                   @r�q��?             @������������������������       �                     @�      �                   (@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   �?���(\��?             $@�      �                   ̅@      �?             @������������������������       �                     �?������������������������       �                     @�      �                   @�8��8��?             @������������������������       �                      @�      �      
            �2@      �?             @������������������������       �                      @�      �                   b�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�                          �?���J�?             6@�      �                   3@�q�q�?             (@�      �                   (@؇���X�?             @������������������������       �                     @������������������������       �                     �?�      �                   �?���Q��?             @������������������������       �                     @������������������������       �                      @                         .@ffffff�?             $@������������������������       �                     @                         �?�$I�$I�?             @������������������������       �                      @                         �?{�G�z�?             @������������������������       �                      @                         @�q�q�?             @������������������������       �                      @������������������������       �                     �?
                         @r�q��?             @������������������������       �                     @������������������������       �                     �?      |                   @�y�����?�            @p@      )                   4�@��-hL��?u            �f@      "                   0�@     ��?             @@                         �?r�q��?             8@            
             %@      �?             @������������������������       �                     @������������������������       �                     �?      !      	            v�@�(\����?             4@                         @ףp=
��?             $@                         B@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         @0�����?             @                         �?z�G�z�?             @������������������������       �                     @                      @33�?      �?              @������������������������       �                     �?������������������������       �                     �?             
             $@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@#      (                   &@      �?              @$      '                   '@؇���X�?             @%      &      
             "@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?*      c                   +@��K�G�?]            �b@+      b                  �O@�ʅʿ��?L            @_@,      ;      	            N�@��63���?J            @^@-      2      	            4�@*
;&���?             G@.      1                ����?`2U0*��?             9@/      0                   �?�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@������������������������       �        	             ,@3      :                  @F@����X�?             5@4      7      
             @�eP*L��?             &@5      6                   d�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @8      9                   �?�q�q�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     $@<      W                ��� @{��;��?+            �R@=      P                ����?�����?            �H@>      O      	            h�@�g�m��?            �B@?      H                   <@����]}�?             ;@@      E                   @*x9/��?             ,@A      B                   �?�<ݚ�?             "@������������������������       �                     @C      D      	            �@      �?             @������������������������       �                      @������������������������       �                      @F      G                   @���Q��?             @������������������������       �                     @������������������������       �                      @I      J      
             %@8�Z$���?             *@������������������������       �                      @K      L                   �?���Q��?             @������������������������       �                      @M      N                  �C@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@Q      V                   ��@r�q��?             (@R      S                   ��@�C��2(�?             &@������������������������       �                      @T      U                  �6@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?X      _                  @G@y0��k��?             :@Y      ^      	            9�@*D>��?	             *@Z      [                   �?r�q��?             @������������������������       �                     @\      ]                pff@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @`      a      	            �@�θ�?             *@������������������������       �                     $@������������������������       �                     @������������������������       �                     @d      k                   @�q�q�?             8@e      j                   @����S�?             ,@f      g                   �?VUUUUU�?             @������������������������       �                     �?h      i                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@l      o                   �?ףp=
��?	             $@m      n                   @      �?              @������������������������       �                     �?������������������������       �                     �?p      w                   @      �?              @q      v                  �1@z�G�z�?             @r      s                   �@�q�q�?             @������������������������       �                     �?t      u                  @K@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @x      y                  �0@�q�q�?             @������������������������       �                     �?z      {                   �?      �?              @������������������������       �                     �?������������������������       �                     �?}      �      	            R�@;C9�v�?2            �S@~      �                  �>@
�N� ��?            �A@      �                   �@ 9�����?             6@�      �                `ff @���Q��?             .@�      �      	            ڐ@�eP*L��?             &@������������������������       �                     @������������������������       �                     @������������������������       �                     @�      �                  �3@և���X�?             @������������������������       �                      @�      �      
             )@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �      
            �3@*D>��?	             *@�      �                   @�g���e�?             &@�      �                `ff�?      �?              @�      �      	            Җ@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                      @�      �                   '@�Ra����?             F@�      �                   @`2U0*��?             9@�      �                  �0@r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �        
             3@�      �      
             @���y4F�?             3@�      �                   ;@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                   1@@4և���?             ,@�      �                   #@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�t�b��%     h�h(h+K ��h-��R�(KM�KK��hb�B t       �z@     0x@     Pz@     �v@      V@      Y@      \@      W@     �M@      T@     �R@     @Q@      *@      :@      @      (@      *@      :@      @              @      @      �?              �?      @      �?              �?              �?                              �?              �?                                      @                      @                              @      6@      @              @                              @      6@      @              �?      4@       @                      �?       @                               @                      �?                      �?      3@                              (@                      �?      @                      �?      �?                      �?                                      �?                              @                       @       @      �?                       @      �?                       @                                      �?               @                                              @      (@                      �?      (@                      �?      @                              @                      �?                                      "@                       @              G@      K@     �P@     �L@     �E@      @@     �O@     �I@      (@       @      (@      @      @       @       @              @               @              @              �?                              �?              @                                              �?               @       @                              �?                       @      �?                       @                                      �?                      @              $@      @      @                                              $@      @                      @                              @      @                       @                               @      @                       @                                      @      ?@      >@     �I@      H@      �?      @       @      &@              @                      �?       @       @      &@      �?       @       @      @               @       @      �?                       @      �?                       @                                      �?               @                      �?                      @                              @      �?                                                      @      >@      9@     �H@     �B@      6@      &@      0@      2@      6@      "@      "@      ,@      5@      �?                      @      �?                      @                                      �?                      0@                              �?       @      "@      ,@                       @              �?       @      �?      ,@      �?       @      �?                       @      �?                      @                              @      �?                      @                                      �?              �?                                                      ,@               @      @      @                      @                       @      �?      @              �?              @              �?                                              @              �?      �?                              �?                      �?                       @      ,@     �@@      3@       @      ,@      6@      2@       @      ,@      @              @       @      @              �?              @              �?                                              @              @       @                               @                      @                               @      (@      �?                              �?               @      (@                       @                                      (@                                      0@      2@                      @      �?                      @                                      �?                      $@      1@                      @                              @      1@                      @                               @      1@                       @      @                       @                                      @                              *@                      &@      �?                      $@                              �?      �?                              �?                      �?              @      6@      @      @      �?      "@      @      @                              @      �?      "@      @                       @                      �?      �?      @              �?              @              �?               @                               @              �?                                              �?                      �?                       @      *@      �?      �?               @                       @      @      �?      �?      �?      @              �?      �?                                      @              �?              @                                              �?      �?              �?              �?                                              �?              =@      4@      C@      7@      <@      ,@     �B@      5@      0@      @      "@      "@                       @              0@      @      @      "@      0@       @      @      @      @       @      @      �?                      @              @       @              �?              �?              �?              �?                                              �?      @      �?                              �?                      @                              "@                       @      �?                       @      �?                                                       @       @                                      �?      �?      @              �?      �?       @                               @              �?      �?                      �?                                      �?                                      @      (@      &@      <@      (@              @      @      @              @              @              @                                              @               @      @      �?               @              �?              �?                              �?              �?                              �?              �?                                      @              (@      @      7@       @      @       @      &@              @       @      @              @                                       @      @                       @                                      @                              @              @       @      (@       @      @       @      &@                       @      &@                      �?      &@                              &@                      �?                              �?                      @                                              �?       @                      �?                                       @      �?      @      �?       @      �?      @              �?      �?      �?              �?      �?                                      �?              �?              �?                                              �?              @                                      �?      �?                      �?                                      �?     pu@     �q@     Ps@     �p@     �f@     `b@      e@     @]@      `@      U@     �X@      H@     @\@      U@     �V@      H@     �C@     �B@      0@      ,@      :@     �B@      .@      (@      @              @       @       @              @       @       @                                              @       @                               @                      @              @                              5@     �B@       @      $@      3@     �@@      @      @      0@                              @     �@@      @      @              @      �?      @                               @              @      �?      @              @      �?                      @                                      �?                                      @      @      ;@      @      �?      @      ;@       @      �?      @      0@       @      �?              ,@              �?              @              �?              �?              �?              �?                                              �?              @                              "@                      @       @       @              @                                       @       @                       @                                       @                      &@                                      �?               @      @      @      @              �?              @                               @              �?               @              �?                                               @       @      @      @                              @               @      @                      �?                              �?      @                      �?                                      @                      *@              �?       @      *@                                              �?       @                      �?                                       @     �R@     �G@     �R@      A@     �Q@     �G@     �R@      ?@     �H@      ?@     �A@      5@      ,@      ,@      7@       @              �?      @                      �?                                      @              ,@      *@      1@       @      *@                              �?      *@      1@       @      �?              "@                              @              �?              @              �?                                              @                      *@       @       @              @              �?                              �?              @                              @       @      �?              �?      @                      �?      @                      �?      �?                      �?                                      �?                              @                              �?                      @      @      �?              @              �?                              �?              @                                      @             �A@      1@      (@      3@      4@      0@      (@      0@      @       @       @      �?      @              �?              @                                              �?              @       @      �?      �?              @      �?      �?              @                                      �?      �?                              �?                      �?              @       @                      @      �?                              �?                      @                                      �?                      *@       @      $@      .@                      �?      &@                              "@                      �?       @                      �?                                       @      *@       @      "@      @      @      �?      @       @                      @              @      �?      @       @       @               @      �?       @                      �?       @                                                      �?                       @              @      �?      �?      �?      @                                      �?      �?      �?              �?                                      �?      �?                      �?                                      �?       @      @      @       @      @              �?       @      @                       @                               @      @                              @              �?                              �?              @                              �?      @       @              �?      @      �?                      @      �?                      @                              @      �?                              �?                      @                      �?                                              �?              .@      �?              @      .@                       @      .@                                                       @              �?              �?                              �?              �?                      6@      0@      D@      $@              @      ;@                      @       @                       @       @                       @                                       @                      @                              �?      9@                      �?      $@                              "@                      �?      �?                      �?                                      �?                              .@              6@      $@      *@      $@      0@      "@      *@      $@      .@                              �?      "@      *@      $@      �?      @      @      $@               @      @      $@              �?       @       @              �?       @       @                       @      �?                       @                                      �?              �?              �?                              �?              �?                                              @              �?       @       @                               @              �?       @                      �?                                       @              �?      @                              @                      �?                                      @      "@                              @                      @      @                      @      �?                      �?      �?                              �?                      �?                              @                                      @              @      �?                              �?                      @                              @                      @       @                              �?                      @                               @      �?                      �?      �?                                                      �?      0@              @              0@                                              @             �J@     �O@     �Q@     @Q@      F@      =@     �C@      7@      B@      ,@      3@      &@      5@      *@      0@      $@      0@       @      @      @      �?      �?              @      �?      �?                      �?                                      �?                                              @      .@      @      @       @      .@       @                      @                              "@       @                      "@                                       @                              @      @       @              @      �?      �?                      �?                      @              �?              @                              �?              �?                              �?              �?                                      @      �?                              �?                      @              @      @      (@      @      �?      @      &@      �?      �?      @      @      �?              @              �?              �?              �?                              �?              �?                              @                      �?              @                              @              �?                                              @              @      �?      �?       @              �?      �?       @              �?               @              �?                                               @                      �?              @                              .@      �?      @      �?      �?      �?       @      �?      �?      �?              �?              �?                      �?                      �?                              �?      �?                                               @              ,@              �?                              �?              ,@                               @      .@      4@      (@       @      .@      �?               @      *@      �?                      *@      �?                      �?      �?                              �?                      �?                              (@                       @                              @       @                              �?                      @      �?                      @                                      �?                                      3@      (@                      3@      @                      3@      �?                      "@      �?                       @                              �?      �?                      �?                                      �?                      $@                                      @                              @      "@      A@      @@      G@      �?      @              3@                              "@      �?      @              $@              @              @              @               @               @                               @               @               @                                               @                              @      �?       @              @      �?      �?                      �?                                      �?                              �?              @              �?              �?              �?                                              �?                              @       @      <@      @@      ;@       @      6@      .@      @       @      6@      @              �?      @      @              �?      @      @              �?      @                      �?                                      @                                      @                       @                      �?      .@      �?                              �?              �?      .@                      �?                                      .@                                       @      @                      �?      @                      �?                                      @                      @       @                              �?                      @      �?                      @                               @      �?                              �?                       @              @      @      1@      5@      �?      @      �?                      @                      �?              �?              �?                                              �?              @       @      0@      5@      �?      �?      @      1@      �?                       @                               @      �?                                      �?      @      .@                      @      @                      @      �?                      �?      �?                              �?                      �?                              @                                      @              �?              "@                              "@              �?                      @      �?      &@      @      @      �?      @      @      @      �?      @      �?      @                                      �?      @      �?              �?                                      @      �?                              �?                      @                              �?      @                      �?      �?                      �?                                      �?                               @                      @              d@     �a@     �a@      c@      =@      @      @      �?      =@      �?      @      �?      =@                                      �?      @      �?                      @      �?                              �?                      @                      �?                              @                     �`@     �`@      a@     �b@     @Q@     @P@      V@     @R@      I@     �F@      E@      K@      2@      >@      B@      <@              "@      @      @               @               @              @                              @               @               @               @                               @               @                               @                              �?      @      @              �?              @              �?                                              @                      @      �?                      @                                      �?      2@      5@     �@@      5@              @      @                      �?      @                      �?                                      @                      @                      2@      .@      >@      5@      2@      *@                      (@      �?                      (@                                      �?                      @      (@                              @                      @      @                      @      �?                       @      �?                       @                                      �?                      @                                      @                               @      >@      5@                      @      2@                      @      2@                      @                                      2@                      @                       @      7@      @               @      0@      @               @                                      0@      @                      @      @                      @                                      @                      "@                              @              @@      .@      @      :@      2@      �?              "@      "@                      @                              @      "@                       @      "@                                                       @      "@      �?              @      "@                                      �?              @              �?                                              @      ,@      ,@      @      1@      ,@      ,@      @              "@      @                      "@                                      @                      @      &@      @              @       @                      @                                       @                              @      @                      @                                      @                               @      1@                       @      @                       @      �?                      �?                              �?      �?                              �?                      �?                                       @                              ,@      3@      4@      G@      3@       @      @      *@      @       @      @      (@              �?      @      (@              �?      @      @                              @              �?      @                      �?      �?                              �?                      �?                                       @                                       @              �?      @                              @                      �?                                              �?      @                              @                      �?              1@      ,@     �@@      *@      @      @      @      @      @              @       @      @                                              @       @                              �?                      @      �?                              �?                      @              @      @              @      @       @              @      @                                       @              @               @                                              @              @                      &@      @      ;@       @      &@      @      6@       @                      @              &@      @      .@       @       @      @      @      �?      @      @      @      �?      �?              @                              @              �?               @                               @              �?                              @      @              �?      @      �?                              �?                      @                               @      @              �?       @                                      @              �?               @                              �?              �?              �?                                              �?       @                              @       @      $@      @              �?       @      @              �?      @                              @                      �?                                       @      @                              @                       @              @      �?       @      @      @                                      �?       @      @                               @              �?       @       @                       @                      �?               @                               @              �?                              �?      @                              @                      �?                     �O@     �Q@     �H@     �S@      I@      L@      B@     �C@      @      @      &@      &@      @      @      @      $@      @      �?                      @                                      �?                       @      @      @      $@       @      @      @              �?       @                      �?                                       @                      �?      �?      @                      �?      @                              @                      �?      �?                      �?                                      �?              �?              �?                              �?              �?                                                      $@      �?              @      �?                      @      �?                       @      �?                              �?                       @                              @              �?                              F@      J@      9@      <@     �D@     �A@      9@      8@     �D@      ?@      9@      8@     �C@      @                      8@      �?                      $@      �?                              �?                      $@                              ,@                              .@      @                      @      @                      �?      @                      �?                                      @                      @       @                      @                                       @                      $@                               @      8@      9@      8@       @      "@      8@      ,@       @      "@      ,@      (@       @      "@      ,@       @       @      "@      @               @      @                              @                       @       @                       @                                       @                               @      @                              @                       @                                      &@       @                       @                              @       @                       @                              �?       @                      �?                                       @                              $@                      $@       @                      $@      �?                       @                               @      �?                       @                                      �?                              �?              .@      �?      $@              @      �?      @              @      �?                      @                              �?      �?                              �?                      �?                                              @              $@              @              $@                                              @              @                      @      1@              @      �?      (@              �?      �?      �?              �?      �?                                      �?              �?                              �?              �?                              &@                       @      @              @      �?                      �?                              �?      �?                              �?      @               @      �?      @                      �?       @                              �?                      �?      �?                      �?                                      �?                               @                              �?               @                              �?              �?              �?              �?                                              �?      *@      ,@      *@     �C@      *@      ,@       @              @      *@      @              @      "@                      @      @                      @                                      @                              @                              @      @                               @                      @      �?                              �?                      @                      @      �?      @              @      �?      @              @      �?      @                      �?      @                      �?                                      @              @                              @                                               @                              @     �C@                      �?      8@                      �?      @                      �?                                      @                              3@                      @      .@                      @       @                      @                                       @                      �?      *@                      �?      @                              @                      �?                                      $@�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJC�NhG        hNhG        hHKhIKhJh(h+K ��h-��R�(KK��hb�C               �?       @      @�t�bhVhghQC       ���R�hkKhlhoKh(h+K ��h-��R�(KK��hQ�C       �t�bK��R�}�(hKhyM'hzh(h+K ��h-��R�(KM'��h��B��         4       
             @�+e���?�            �@                           "�@�G�z��?5             T@                           p�@8�#�(�?            �@@                        ���@X�<ݚ�?             "@              	            ��@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @	                            @�q�q�?             8@
                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?                           �?b>���?             5@                           �?$�q-�?             *@                           @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@                           �?      �?              @                           @�q�q�?             @������������������������       �                      @������������������������       �                     �?                           X�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @       /       	            �@})Z6K�?             �G@       $                    �?���%&�?            �B@       !                    @�&5D�?
             1@                            @      �?              @                           �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @"       #       	            �@�����H�?             "@������������������������       �                     �?������������������������       �                      @%       *                    �?�Q����?             4@&       '                    @����X�?	             ,@������������������������       �                     @(       )                    Ι@      �?              @������������������������       �                     @������������������������       �                     @+       ,                    �?�q�q�?             @������������������������       �                     @-       .                 @33�?�q�q�?             @������������������������       �                      @������������������������       �                     �?0       3                    �?ףp=
�?	             $@1       2       	            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @5                       033�?�H�O���?�           ��@6       I                    @JQ8����?           P|@7       <       
             @����bo�?            �A@8       9                    @      �?              @������������������������       �                     @:       ;       	            $�@���Q��?             @������������������������       �                     @������������������������       �                      @=       >       	            ��@|	�%���?             ;@������������������������       �                     @?       F                    %@      �?             8@@       E                    Z�@AA�?             5@A       B                    �?j�V���?             &@������������������������       �                      @C       D                    ��@�����H�?             "@������������������������       �                      @������������������������       �                     �?������������������������       �                     $@G       H       	            n�@�q�q�?             @������������������������       �                     �?������������������������       �                      @J       �       	            �@���O��?
            z@K       �                    )@�׫��?�            �p@L       k                    �?R�bT���?�            �n@M       T       	            ؐ@D^�����?+            �P@N       S                    @ ��WV�?             :@O       P                    �?z�G�z�?             @������������������������       �                     @Q       R                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     5@U       f                    ��@R���Q�?             D@V       ]                    �@�f>����?             =@W       X                    @     ��?             0@������������������������       �                     "@Y       Z                    �?:/����?             @������������������������       �                     @[       \                   �@@      �?             @������������������������       �                      @������������������������       �                      @^       c                    @޾�z�<�?
             *@_       b       	            Ι@��!pc�?             &@`       a                   �=@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@d       e                    �?      �?              @������������������������       �                     �?������������������������       �                     �?g       h       
             %@�C��2(�?             &@������������������������       �                     @i       j                    &@z�G�z�?             @������������������������       �                     �?������������������������       �                     @l       �                    �?��a���?p            `f@m       x       	            ��@���k�?6             W@n       q                    �?8�Z$���?            �C@o       p                    ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @r       w                    @�����H�?             B@s       t                    $�@�<ݚ�?             2@������������������������       �        	             *@u       v                    *@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     2@y       �       
             !@��]ۡ�?            �J@z       �                    K@������?             ,@{       �                    ��@�Q����?             $@|       }                    @      �?              @������������������������       �                     �?~       �                 ����?؇���X�?             @       �                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                    !@�q�q�?            �C@�       �                    "�@���Q��?             @������������������������       �                     @������������������������       �                      @�       �                    $@��)��?             A@�       �                    �?     ��?             @@������������������������       �                     �?�       �                    @���M�?             ?@�       �                 ����?�C��2(�?             6@������������������������       �                     ,@�       �       
             )@      �?              @������������������������       �                     @�       �                    @      �?             @������������������������       �                      @������������������������       �                      @�       �                    �@�q�q�?             "@������������������������       �                     @�       �       	            Ɩ@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    @��>x�?:            �U@�       �                    ��@��wC���?-            �P@�       �                    x�@��.k���?             A@�       �                    �?�n_Y�K�?             :@�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @�LQ�1	�?             7@������������������������       �                      @�       �                    %@��S���?	             .@�       �       
             /@�<ݚ�?             "@������������������������       �                     @�       �                    ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                 ����?r�q��?             @�       �                    .@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @�       �                    @     ��?             @@�       �       
             /@�5�;N��?             9@�       �                   �2@�E�_���?             5@�       �       	            {�@�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?�       �                   �;@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @      �?             @������������������������       �                     �?�       �                    @�q�q�?             @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    �?և���X�?             @������������������������       �                      @�       �                    ��@���Q��?             @������������������������       �                     �?�       �                    ��@      �?             @������������������������       �                      @�       �       	            �@      �?              @������������������������       �                     �?������������������������       �                     �?�       �       
             1@����X�?             5@�       �       	            Ζ@���y4F�?             3@������������������������       �        	             .@������������������������       �                     @������������������������       �                      @�       �                    $@(������?             3@������������������������       �                     �?�       �       	            h�@�)O�?
             2@�       �                    ��@�8��8��?             @�       �                    �?�q�q�?             @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     (@�       	                  @K@�����?d            @c@�             
            �1@����C�?V            ``@�       �       
             @�)S;��?K            �[@�       �       	            ݨ@">�֕�?            �A@�       �                    t�@8�Z$���?	             *@������������������������       �                     $@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     6@�       �                    @"!h�3��?5            �R@�       �                    ?@r�q��?             8@�       �                    H�@��\���?             1@�       �                    �?H�z�G�?             $@�       �                    ܂@������?             @�       �                    �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @������������������������       �                     @�       �                    ֗@;h����?"            �I@�       �       	            ݪ@L�߮V�?            �C@�       �       	            �@�m펠�?            �@@�       �                    @j�V���?             &@�       �                    �?      �?             @������������������������       �                     �?�       �                    ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     6@�       �                    �?      �?             @������������������������       �                      @�       �                   �>@      �?             @������������������������       �                     �?������������������������       �                     @�                          @r�q��?             (@�                           %@�����H�?             "@������������������������       �                      @������������������������       �                     �?            	            (�@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         ,�@&%�ݒ��?             5@                         �@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �        	             1@
            	            �@�p�F�:�?             7@������������������������       �                      @                        �O@AA�?             5@            
             /@�IєX�?             1@������������������������       �                     &@                         �?r�q��?             @                         @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                         @      �?             @������������������������       �                      @������������������������       �                      @      >                   �@�Rq<��?�           ��@      ;                   @a�O���?h           ȁ@      :                   ��@}��7�?6             V@      9                    �@�c�i���?3            @T@      "      	            ʞ@&�(f���?0            @S@            	            6�@$�q-�?            �C@������������������������       �                    �@@                         @      �?             @������������������������       �                      @       !                  �D@      �?             @������������������������       �                     @������������������������       �                     �?#      2      	            ��@�p9W���?             C@$      '                   �?�\��N��?             3@%      &      	            Ȣ@r�q��?             @������������������������       �                     �?������������������������       �                     @(      )                  �8@*D>��?	             *@������������������������       �                     �?*      +                   ��@�q�q�?             (@������������������������       �                     @,      1                   ��@�<ݚ�?             "@-      0                   t�@���Q��?             @.      /                ���@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @3      8                `ff @�KM�]�?             3@4      7                   �@      �?              @5      6                   �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     &@������������������������       �                     @������������������������       �                     @<      �                `ff @��&c��?2           ~@=      �                   �?38@)��?�            pq@>      o                   +@�ۦ�qA�?o             f@?      l                   ~�@���X�??            �X@@      E                   �?�C4T2�?;             W@A      B      	            8�@�q�q�?             5@������������������������       �        	             .@C      D                   �?�q�q�?             @������������������������       �                      @������������������������       �                     @F      Y                   ��@�ߌJ���?.            �Q@G      V                   @�کB���?             =@H      I                   .@����Gc�?             3@������������������������       �                     @J      U                   L@�q-��?             *@K      T                   #@��ˠ�?	             &@L      S                   �?      �?              @M      N                   @�8��8��?             @������������������������       �                     �?O      R                ����?�Q����?             @P      Q      	            >�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     @������������������������       �                      @W      X      	            ��@�z�G��?             $@������������������������       �                     @������������������������       �                     @Z      k      	            Ӧ@$I�$I��?             E@[      d                   �?�'s�	U�?             A@\      ]                   �?>;n,��?             &@������������������������       �                     @^      a                   @      �?              @_      `      	            �@�q�q�?             @������������������������       �                      @������������������������       �                     �?b      c                033�?z�G�z�?             @������������������������       �                     @������������������������       �                     �?e      f                   @D%��N��?             7@������������������������       �                     @g      j                   @�IєX�?	             1@h      i                ����?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@������������������������       �                      @m      n      
             @r�q��?             @������������������������       �                     �?������������������������       �                     @p      �                   �?puqrZC�?0            �S@q      z                   �?�^)��?             9@r      s                  @B@hE#߼�?             .@������������������������       �                     "@t      u                   �?�8��8��?             @������������������������       �                     �?v      w      
             $@{�G�z�?             @������������������������       �                      @x      y      	            ,�@�q�q�?             @������������������������       �                      @������������������������       �                     �?{      |                   @���(\��?             $@������������������������       �                     @}      ~                   �?      �?             @������������������������       �                     �?      �      
             @z�G�z�?             @������������������������       �                      @�      �                   6@�q�q�?             @������������������������       �                     �?�      �                  �0@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   @��;F��?              K@�      �      	            �@�˹�m��?             3@������������������������       �                     $@�      �      	            ��@��E���?             "@�      �      
             /@r�q��?             @������������������������       �                     @������������������������       �                     �?�      �                   ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �      	            7�@
�N� ��?            �A@�      �                ����?3������?             =@�      �      
             @     @�?             0@�      �                ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   &@
ц�s�?
             *@�      �      	            ��@H�z�G�?             $@������������������������       �                     @�      �      
             /@؇���X�?             @������������������������       �                     @�      �      	            ՠ@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   0@8�Z$���?             *@�      �                   |�@���Q��?             @������������������������       �                     �?�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                  @N@"h��:��?F            �Y@�      �                   '@UC����?B            �W@�      �                   �?�-P��?7            @S@�      �                033�?     P�?             @@�      �                   @n����?             =@������������������������       �                     @�      �      
             '@�"AM�h�?             :@�      �      
             #@      �?
             (@�      �                  �;@VUUUUU�?             "@�      �      	            ��@���Q��?             @������������������������       �                      @������������������������       �                     @�      �      	            ��@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �      	            F�@/����?             ,@������������������������       �                     @�      �      	            _�@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?�      �                   ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   0�@|6)���?             �F@�      �                    @*�c{��?             3@�      �                   �?0�����?             @�      �                   �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �      
             @�q�q�?             (@������������������������       �                      @�      �      	            š@��(\���?             $@�      �                033�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                   '@G���ջ�?             :@�      �                   �?     ��?             0@�      �                  �L@և���X�?             @�      �                   @���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @������������������������       �                     "@�      �                   @{�G�z�?             $@�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @�      �                   �?      �?             @������������������������       �                     �?�      �                   @z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �      	            ��@=[y���?             1@�      �      
             1@����X�?             @������������������������       �                     @������������������������       �                      @�      �                   :@ףp=
�?             $@�      �      	            �@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @�                         +@Pϳ;=8�?}            @i@�      
      
             !@�ٴ��?F             [@�      �                   �?VUUUU�?              H@�      �                  �5@s
^N���?             <@�      �                   �?>4և���?             ,@�      �      
             @B{	�%��?             "@������������������������       �                     �?�      �                   @      �?              @������������������������       �                     @������������������������       �                     �?�      �                   %@���Q��?             @������������������������       �                      @������������������������       �                     @�      �      	            �@�X�C�?
             ,@�      �                   �?�����H�?             "@�      �      	            �@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                   @���Q��?             @������������������������       �                      @������������������������       �                     @�                         %@�G�z��?             4@�                         @���Er�?             1@                          �?�m۶m��?             ,@������������������������       �                     �?            	            @.y0��k�?             *@������������������������       �                     &@                         ԉ@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @      	                  �E@�q�q�?             @������������������������       �                     �?������������������������       �                      @                         ؃@�������?&             N@                         @ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@            	            ��@��h o��?!             I@������������������������       �                     3@            	            ʩ@w���<�?             ?@            	            �@�C��2(�?             6@            	            ��@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     2@                         @�<ݚ�?             "@                         @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @      /                   ��@$g�P��?7            �W@      "      	            ��@�j����?&            @Q@      !                   -@h�����?             <@                       ���@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     7@#      (      	            $�@���e��?            �D@$      %      	            m�@z�G�z�?	             4@������������������������       �                     &@&      '                  �G@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @)      .                   �@؇���X�?             5@*      +                   @      �?              @������������������������       �                     @,      -                   @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     *@0      3                   @��d�`T�?             9@1      2      	            @z�G�z�?             @������������������������       �                     �?������������������������       �                     @4      7                   ,@>
ףp=�?             4@5      6      
             /@      �?              @������������������������       �                     �?������������������������       �                     �?8      ;                   �?�ӭ�a��?             2@9      :      	            �@����X�?             @������������������������       �                      @������������������������       �                     @<      =                   @�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@?      �      
            �1@F�u�l}�?5            @@      �      	            U�@~,��}�?           �y@A      �                  �0@x�[�&��?�            �q@B      �                   @w���%��?�            `l@C      b                   �?�
F%u�?C             Y@D      K      	            ��@HPS!���?$             J@E      J                   @���7�?             6@F      G      	            (�@ףp=
�?             $@������������������������       �                      @H      I                   ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@L      _                   @	���ĳ�?             >@M      N                   �?~e�.y0�?             :@������������������������       �                      @O      R                   �?�q�q�?             8@P      Q      	            ��@�����H�?             "@������������������������       �                      @������������������������       �                     �?S      T      
             @�Q����?             .@������������������������       �                      @U      ^                   K@�؉�؉�?
             *@V      [                   ��@��!pc�?	             &@W      Z                   �?�����H�?             "@X      Y                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @\      ]      
             +@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @`      a                  �5@      �?             @������������������������       �                     �?������������������������       �                     @c      �                   @�8��8N�?             H@d      m                   �?b�h�d.�?            �A@e      h                ����?����X�?	             ,@f      g      	            ��@؇���X�?             @������������������������       �                     �?������������������������       �                     @i      l                   @և���X�?             @j      k                   ��@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @n      �                   @ܤ�[r�?             5@o      r                   @�$�_�?             3@p      q                   �?      �?             @������������������������       �                     @������������������������       �                     �?s      t                   @�Q����?	             .@������������������������       �                      @u      ~      
             /@*D>��?             *@v      w                   �?      �?              @������������������������       �                     @x      }                  @M@�Q����?             @y      z                   �?VUUUUU�?             @������������������������       �                     �?{      |      
             @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @      �                   N�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                   �?&�q-�?	             *@�      �      
             !@0�����?             @������������������������       �                     @�      �      	            �@      �?             @������������������������       �                     �?�      �      
             (@�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   @r�q��?             @������������������������       �                     @������������������������       �                     �?�      �                   P�@�(��i��?J            �_@�      �                033@��|��?(             Q@�      �      
            �0@2�[��?            �@@�      �      
             -@     ��?             @@�      �      	            ��@^�`���?             :@�      �                  �6@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @�      �                   -@8߄*�u�?
             1@������������������������       �                     �?�      �                   �?      �?	             0@������������������������       �                     .@������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�      �      	            �@?B+)�9�?            �A@�      �                   �?P���Q�?             4@������������������������       �                     &@�      �                   �?�����H�?             "@�      �                @33@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �      
             #@��S���?             .@������������������������       �                     @�      �                   �@z�G�z�?             $@������������������������       �                      @������������������������       �                      @�      �      	            T�@�Oi�>��?"            �M@�      �                   �?d}h���?             ,@�      �                   &�@      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                      @�      �                   �@(�Q_�?            �F@�      �                   @�8��8��?             8@������������������������       �                     @�      �                   �?p=
ףp�?             4@�      �                ����?      �?              @�      �                   �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @�      �                   ؙ@r�q��?             (@������������������������       �                     �?�      �      	            5�@�C��2(�?             &@������������������������       �                     @�      �      	            ��@z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �                   @�����?             5@�      �      
            �0@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     (@�      �                `ff@�:m���?'             N@�      �                ���@�8��8��?             H@�      �      	            ��@�ƄIUX�?            �E@�      �      
             )@�#*�6�?             ;@�      �                   �?��S�ۿ?             .@�      �                    @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     &@�      �      	            ��@�q�q�?             (@������������������������       �                     @�      �                   �?�����H�?             "@������������������������       �                     @�      �                   @r�q��?             @������������������������       �                     @�      �                   !@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     0@�      �                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @�      �      
             '@�������?             (@�      �                   �?VUUUUU�?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �      	            ؚ@�����H�?             "@������������������������       �                      @������������������������       �                     �?�      �                   ֞@�â��,�?M             _@�      �                   #@��d��?K             ^@������������������������       �        E            �\@�      �                   ,@r�q��?             @������������������������       �                     �?������������������������       �                     @�      �                   +@      �?             @������������������������       �                      @������������������������       �                      @�                         @@]�{��?4            �U@�      �                033@�5��P^�?             C@�      �                   F@*�c{��?             3@�      �                   @@���!pc�?             &@�      �                   @և���X�?             @������������������������       �                      @�      �                   �?���Q��?             @������������������������       �                      @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                   �?      �?              @������������������������       �                     @�      �      
            �2@{�G�z�?             @������������������������       �                      @�      �                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?             	            �@�lO���?	             3@������������������������       �                      @                         8�@�IєX�?             1@������������������������       �                     "@            	            A�@      �?              @������������������������       �                     @������������������������       �                     �?                         +@�t�*�?            �H@                      ����?     ��?             @@	      
                   F@z�G�z�?             @������������������������       �                     �?������������������������       �                     @                         �?VUUUUU�?             ;@                         @*�c{��?	             3@            	            f�@޾�z�<�?             *@                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@                         �?�8��8��?             @                      `ff�?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @            
            �2@      �?              @������������������������       �                      @                         ^�@      �?             @������������������������       �                     @������������������������       �                     @      $                   �?ҳ�wY;�?             1@                      ���@�C��2(�?             &@������������������������       �                     @       #                033@      �?             @!      "                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @%      &      	            ԣ@r�q��?             @������������������������       �                     @������������������������       �                     �?�t�b��J     h�h(h+K ��h-��R�(KM'KK��hb�B�d       �z@     px@     `x@     �x@      1@      4@      @@      &@      $@      @      2@       @      @      �?       @              @      �?                      @                                      �?                                       @              @       @      0@       @       @      �?                       @                                      �?                       @      �?      0@       @                      (@      �?                       @      �?                              �?                       @                              $@               @      �?      @      �?       @      �?                       @                                      �?                                      @      �?                              �?                      @              @      1@      ,@      "@      @      1@      *@              @      @      "@               @      @      �?               @              �?               @                                              �?                      @                      �?               @              �?                                               @              @      (@      @                      $@      @                      @                              @      @                              @                      @                      @       @                      @                              �?       @                               @                      �?                                              �?      "@                      �?      �?                      �?                                      �?                               @     �y@     0w@     `v@     �w@     @]@     @a@     @Z@     @W@      @      @      4@      @      @      @       @                      @                      @               @              @                                               @              @      @      2@      @      @                                      @      2@      @               @      2@      �?               @       @      �?               @                                       @      �?                       @                                      �?                      $@                      �?               @              �?                                               @     �[@     �`@     @U@     �V@     �[@      _@      =@             @[@     �[@      :@              <@      8@      ,@              9@      �?                      @      �?                      @                              �?      �?                      �?                                      �?                      5@                              @      7@      ,@              @      *@      *@               @      &@      @                      "@                       @       @      @                              @               @       @                       @                                       @                      �?       @      $@              �?      �?      "@              �?      �?                              �?                      �?                                              "@                      �?      �?                      �?                                      �?                      $@      �?                      @                              @      �?                              �?                      @                     @T@     �U@      (@             �F@      D@      @             �@@      @                      �?       @                      �?                                       @                      @@      @                      ,@      @                      *@                              �?      @                              @                      �?                              2@                              (@      A@      @              @      @       @              @       @       @              @       @                              �?                      @      �?                      @      �?                              �?                      @                              @                                               @                      @                      @      <@      @              @       @                      @                                       @                      @      :@      @              @      :@      @              �?                               @      :@      @               @      4@                              ,@                       @      @                              @                       @       @                       @                                       @                              @      @                      @                              �?      @                      �?                                      @                               @              B@      G@      @              5@      D@      @              2@      0@                      $@      0@                       @      �?                       @                                      �?                       @      .@                               @                       @      @                      @       @                      @                              �?       @                      �?                                       @                      �?      @                      �?      �?                              �?                      �?                                      @                       @                              @      8@      @              @      5@      �?              �?      3@      �?                      2@      �?                      2@                                      �?              �?      �?                      �?                                      �?                       @       @                      �?                              �?       @                              �?                      �?      �?                      �?                                      �?                              @      @                               @                      @       @                              �?                      @      �?                       @                              �?      �?                      �?                                      �?              .@      @                      .@      @                      .@                                      @                               @                       @      ,@      @              �?                              �?      ,@      @              �?       @      @              �?       @                      �?      �?                              �?                      �?                                      �?                                      @                      (@                               @      L@     �V@              @     �J@      R@              @      J@     �K@                      &@      8@                      &@       @                      $@                              �?       @                      �?                                       @                              6@              @     �D@      ?@              �?      @      1@              �?      @      $@              �?      @      @              �?      @      @              �?              @              �?                                              @                      @                              @                                      @                              @               @     �A@      ,@               @     �@@      @               @      >@      �?               @       @      �?               @      �?      �?                              �?               @      �?                       @                                      �?                              @                              6@                              @      @                       @                              �?      @                      �?                                      @                       @      $@                      �?       @                               @                      �?                              �?       @                      �?                                       @              @      �?      1@              @      �?                      @                                      �?                                      1@               @      @      2@                       @                       @      �?      2@                      �?      0@                              &@                      �?      @                      �?      �?                              �?                      �?                                      @               @               @               @                                               @     Pr@      m@     �o@      r@     �h@      `@     �`@     �[@     �E@      "@      ,@      6@      B@      "@      ,@      6@      B@      "@      ,@      2@      B@      @                     �@@                              @      @                               @                      @      �?                      @                                      �?                              @      ,@      2@              @      (@      �?              �?      @                      �?                                      @                      @      @      �?                              �?              @      @                      @                               @      @                       @      @                      �?      @                              @                      �?                              �?                                      @                               @      1@                       @      @                       @       @                               @                       @                                      @                              &@                              @      @                              c@      ^@     �]@     @V@      V@     @T@      J@      M@      N@      K@     �B@      :@      <@     �D@      (@      1@      7@     �D@      &@      1@              .@       @      @              .@                                       @      @                       @                                      @      7@      :@      "@      *@      (@      @      @      @      "@      @              @      @                              @      @              @      @      @              @      @      @               @      @      �?               @                              �?      @      �?              �?              �?              �?              �?                                              �?      @                                       @                                              @               @                      @              @              @                                              @              &@      5@       @       @      &@      5@       @              @      @      �?              @                               @      @      �?               @      �?                       @                                      �?                              @      �?                      @                                      �?              @      0@      �?              @                                      0@      �?                      @      �?                      @                                      �?                      &@                                               @      @              �?                              �?              @                              @@      *@      9@      "@      0@      @      @              &@      @      �?              "@                               @      @      �?                      �?                       @       @      �?                       @                       @              �?               @                                              �?              @      �?      @              @                              �?      �?      @              �?                                      �?      @                               @                      �?       @                              �?                      �?      �?                      �?                                      �?              0@      "@      4@      "@      &@      @       @      �?      $@                              �?      @       @      �?      �?      @                              @                      �?                                               @      �?                       @                                      �?      @      @      2@       @      @      @      2@       @      @      @      @       @                      �?       @                      �?                                       @      @      @      @              @      �?      @              @                                      �?      @                              @                      �?       @                               @                      �?                              @                       @              &@               @              @              �?                              �?              @                              @              �?                                               @                                      @      <@      ;@      .@      @@      <@      ;@      .@      8@      7@      9@      ,@      .@      "@      0@      �?      @      "@      0@              @              @                      "@      *@              @      @      @              @      @      @              @       @      @                       @                                      @                      �?                      @      �?                                                      @      @                              @      $@              �?      @                                      $@              �?              $@                                              �?                      �?       @                               @                      �?              ,@      "@      *@      "@      �?       @      "@      @              �?      �?      @              �?      �?                      �?                                      �?                                      @      �?      �?       @       @                               @      �?      �?       @              �?      �?                      �?                                      �?                                       @              *@      @      @       @      *@      @                      @      @                       @      @                              @                       @                               @                              "@                                      @      @       @              @              �?                              �?              @                              �?      @      �?              �?                                      @      �?                              �?                      @              @       @      �?      "@      @       @                      @                                       @                                      �?      "@                      �?       @                      �?                                       @                              @                               @     @P@     �C@     �P@      ?@      A@      1@     �F@      (@      .@      ,@      ,@      @      @      "@      (@      @      @      �?      "@      �?              �?      @      �?                              �?              �?      @                              @                      �?                      @               @                               @              @                              �?       @      @       @      �?       @                      �?      @                      �?                                      @                              @                                      @       @                               @                      @              &@      @       @       @      &@      @      �?              &@       @      �?                      �?                      &@      �?      �?              &@                                      �?      �?                              �?                      �?                              @                                      �?       @                      �?                                       @      3@      @      ?@      @              �?      "@                      �?                                      "@              3@       @      6@      @      3@                                       @      6@      @               @      4@                       @       @                               @                       @                                      2@                               @      @                       @       @                               @                       @                                      @      ?@      6@      6@      3@      ;@      1@      @      2@      ;@      �?                      @      �?                      @                                      �?                      7@                                      0@      @      2@              0@      @                      &@                              @      @                      @                                      @                              @      2@                      @      @                              @                      @      �?                      @                                      �?                              *@      @      @      .@      �?      �?      @                      �?                                      @                      @      �?      .@      �?      �?      �?                      �?                                      �?                       @              .@      �?       @              @               @                                              @                              $@      �?                              �?                      $@             @X@      Z@      ^@      f@     @T@     �S@      [@     �a@     @T@     �S@     @Z@      6@     �R@      H@     �T@      5@     �D@      ;@      :@      @      5@      2@      @      @      5@      �?                      "@      �?                       @                              �?      �?                      �?                                      �?                      (@                                      1@      @      @              1@      @      @                       @                      1@      @      @               @      �?                       @                                      �?                      "@      @      @                       @                      "@      �?      @              "@      �?      �?               @      �?                      @      �?                              �?                      @                              @                              �?              �?              �?                                              �?                               @                      �?      @                      �?                                      @      4@      "@      3@              ,@      @      2@              @              $@              �?              @              �?                                              @              @              @              @               @              @                                               @                               @              $@      @       @              $@      �?       @              @              �?              @                                              �?              @      �?      @                               @              @      �?      @              @      �?      �?              @                              @      �?      �?              �?      �?      �?              �?                                      �?      �?                              �?                      �?                       @                              �?              @              �?                                              @                       @                      @      @      �?              �?      @      �?                      @                      �?       @      �?              �?                                       @      �?                              �?                       @                      @      �?                      @                                      �?                      A@      5@     �L@      .@      7@      .@      =@      �?      @      @      5@      �?      @      @      5@      �?      @      @      .@      �?      @      @                      @                                      @                              �?      .@      �?                              �?              �?      .@                              .@                      �?                                      @                      �?                      3@       @       @              3@      �?                      &@                               @      �?                      @      �?                      @                                      �?                      @                                      @       @                      @                               @       @                               @                       @                      &@      @      <@      ,@      &@      @                      @      @                              @                      @                               @                                      @      <@      ,@              �?      "@      ,@                              @              �?      "@      $@              �?      @                      �?       @                               @                      �?                                      @                               @      $@                      �?                              �?      $@                              @                      �?      @                      �?                                      @               @      3@                       @      @                              @                       @                                      (@              @      ?@      6@      �?      @      6@      5@              @      6@      1@              @      6@      �?              �?      ,@                      �?      @                              @                      �?                                      &@                      @       @      �?              @                                       @      �?                      @                              @      �?                      @                               @      �?                              �?                       @                                      0@              �?              @              �?                                              @              �?      "@      �?      �?      �?      �?              �?      �?                      �?                              �?      �?                                      �?                               @      �?                       @                                      �?                              @     @^@                      �?     �]@                             �\@                      �?      @                      �?                                      @                       @       @                       @                                       @      0@      9@      (@      A@      @      5@       @      $@      @      @      �?      $@      @                       @      @                      @                               @      @                       @       @                              �?                       @      �?                                                       @                              @              @      �?       @              @                               @      �?       @                               @               @      �?                       @                                      �?               @      0@      �?               @                                      0@      �?                      "@                              @      �?                      @                                      �?              &@      @      $@      8@      &@      @      @      *@      @      �?                              �?                      @                              @      @      @      *@      @      @      �?      $@       @      �?              $@       @      �?                              �?                       @                                                      $@      @       @      �?                       @      �?                              �?                       @                      @                               @              @      @       @                                              @      @                              @                      @                              @      &@                      �?      $@                              @                      �?      @                      �?      �?                      �?                                      �?                               @                      @      �?                      @                                      �?�t�bubhhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�R�[hG        hNhG        hHKhIKhJh(h+K ��h-��R�(KK��hb�C               �?       @      @�t�bhVhghQC       ���R�hkKhlhoKh(h+K ��h-��R�(KK��hQ�C       �t�bK��R�}�(hKhyM�hzh(h+K ��h-��R�(KM���h��Bx�         p                   �?�n����?�            �@       �       	            w�@�bx���?           ��@       0                    �?�d���?           �x@                           �@K���@�?@            �Y@������������������������       �                     "@              	            H�@�5v���?;            �W@                           @�:�]��?            �I@                          �1@��?^�k�?            �A@	       
                    @      �?              @������������������������       �                     @������������������������       �                     �?������������������������       �                     ;@                           ��@     ��?             0@������������������������       �                     (@                           @      �?             @������������������������       �                     @������������������������       �                     �?       #                    @Fc�[���?            �E@                           �?�8��8��?             2@������������������������       �                      @       "                   @E@     ��?             0@                           �?
ц�s�?
             *@              	            �@h/�����?             "@                        ����?����X�?             @������������������������       �                     @                           L�@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @       !                   �=@      �?             @                            �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @$       '       
             @`�Q��?             9@%       &                 ����?      �?              @������������������������       �                     �?������������������������       �                     �?(       )                    @X��t��?             7@������������������������       �                     �?*       /                    �?���7�?             6@+       ,                    �?�8��8��?             (@������������������������       �                     @-       .                 ����?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     $@1       b                    ��@��OD�7�?�            @r@2       7                    �?�ЬS��?Q            �^@3       6                    *@"pc�
�?            �@@4       5       	            F�@     ��?             @@������������������������       �                     ;@������������������������       �                     @������������������������       �                     �?8       U                    +@02�5���?<            �V@9       D                    �?&�X�%�?'             N@:       C                   @@@      �?             @@;       <       
             @E�ϣ1��?             3@������������������������       �                     @=       B                    �?H�7�&��?             .@>       A                    T�@{�G�z�?             @?       @                    �@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     $@������������������������       �                     *@E       P                    x�@���>4��?             <@F       M                    @     ��?             0@G       L                    #@�θ�?	             *@H       K                    @���Q��?             @I       J                   �D@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @N       O                 @33�?�q�q�?             @������������������������       �                     �?������������������������       �                      @Q       R                    @�q�q�?             (@������������������������       �                      @S       T       	            B�@z�G�z�?             $@������������������������       �                      @������������������������       �                      @V       a       
             /@r�q��?             >@W       ^                    �?      �?             4@X       Y                    �?X�<ݚ�?             "@������������������������       �                     @Z       [                   �@@�q�q�?             @������������������������       �                     @\       ]                 ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @_       `                 pff@�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?������������������������       �                     $@c       �                    @�M���?r             e@d       �                    �?�䣓�N�?U            �_@e       ~                 `ff�?��"AM�?$             J@f       w                 ����?��T�	��?             E@g       p                    @���6c�?             A@h       o                    @�M�]��?             1@i       l                    �?8�Z$���?             *@j       k                    ,@r�q��?             @������������������������       �                     �?������������������������       �                     @m       n       	            �@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @q       r                    #@@�0�!��?	             1@������������������������       �                     �?s       t                    �?      �?             0@������������������������       �                     $@u       v       	             �@�q�q�?             @������������������������       �                     @������������������������       �                      @x       y                    @      �?              @������������������������       �                      @z       }       	            �@�8��8��?             @{       |                    2@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @       �                    !@ףp=
�?             $@�       �       
             /@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	            ��@V������?1            �R@�       �       	            ��@r�q��?             2@������������������������       �                     @�       �       
             '@      �?             (@�       �                   �F@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�       �       	            x�@H�$I�$�?%             L@�       �                   @K@г�wY;�?             A@������������������������       �                     ?@�       �                    0@�q�q�?             @������������������������       �                     �?������������������������       �                      @�       �                    �?"pc�
�?             6@�       �                 033�?�q�q�?             @�       �                    @z�G�z�?             @������������������������       �                      @�       �       
             @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?      �?
             0@�       �                    �@�<ݚ�?             "@�       �                    @      �?              @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �       	            �@�҇����?            �E@������������������������       �                     1@�       �                    �?y0��k��?             :@�       �                    ��@.y0��k�?             *@�       �                    �@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                    D�@�	j*D�?
             *@�       �                    @      �?	             (@������������������������       �                      @�       �                    �?      �?             @������������������������       �                     �?�       �                    .�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?�                          @j)�1U��?           pz@�       �                    �?���k��?w            @g@�       �       
             @B������?            �G@�       �                    �?���Q��?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @�       �                    @����>�?             E@�       �       
             %@�ˠT�?            �@@�       �                    �?�����H�?	             2@������������������������       �                     (@�       �                    8@�q�q�?             @������������������������       �                      @������������������������       �                     @�       �                    #@�.�?��?             .@������������������������       �                     �?�       �       	            Х@X�Cc�?             ,@������������������������       �                      @�       �                    �?r�q��?             @������������������������       �                     @�       �       
             .@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�       �                    �?y�s��?[            `a@�       �                    �?C��6�?!             I@�       �                    �?��#��Z�?             6@�       �                 033@      �?             ,@�       �                    @�$I�$I�?             @�       �                   �J@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?      �?              @�       �                    Z�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @z�G�z�?             @������������������������       �                     @������������������������       �                     �?�       �                    @      �?             <@�       �       
             /@ҳ�wY;�?             1@�       �                    ��@�eP*L��?             &@�       �                    ��@r�q��?             @������������������������       �                     �?������������������������       �                     @�       �                   @E@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�       �                    @���!pc�?             &@�       �                    �?���Q��?             @������������������������       �                      @�       �       	            w�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�              
             $@� W<>�?:            @V@�       �                 033@~fL���?            �@@�       �                    (�@�
�[-�?             =@������������������������       �                     "@�       �       	            
�@�Q����?             4@�       �                    C@      �?             @������������������������       �                      @������������������������       �                      @�       �                    L@      �?
             0@������������������������       �                     (@�       �                    @      �?             @������������������������       �                     �?������������������������       �                     @�       �                 pff@      �?             @�       �       	            -�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @                         ��@ܶm۶m�?%             L@                         @UP��g��?             G@                         �?9��8���?             8@������������������������       �                     �?            	            ��@�2'�%�?             7@                         �?      �?             (@������������������������       �                      @                         �?z�G�z�?             $@	      
                   @      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @            	            ��@�C��2(�?             &@������������������������       �                     @            	            L�@r�q��?             @������������������������       �                     �?������������������������       �                     @                         @8�A�0��?             6@������������������������       �                      @                        �A@��X��?
             ,@                      `ff�?      �?              @������������������������       �                     @                         0@�Q����?             @                         @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     $@      c      	            @�@B�QU���?�            �m@      *                  �0@+��K��?]            �b@       #                  �1@     ��?             @@!      "      
            �3@���7�?             6@������������������������       �                     5@������������������������       �                     �?$      )      	            ܧ@���Q��?             $@%      &                   ��@      �?              @������������������������       �                     @'      (                   1@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                      @+      F                   ��@d���5�?J            �]@,      ;                   !@��X���?             �I@-      0                   ��@8߄*�u�?             A@.      /                  �9@�q�q�?             @������������������������       �                      @������������������������       �                     @1      :                  �I@@4և���?             <@2      3                   @�r����?             .@������������������������       �                     "@4      7                   �?�q�q�?             @5      6                   H@      �?             @������������������������       �                     @������������������������       �                     �?8      9                   6@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     *@<      =                  �0@ҳ�wY;�?
             1@������������������������       �                     @>      ?                  @@@�eP*L��?             &@������������������������       �                     @@      A                   �?      �?              @������������������������       �                     �?B      E                   �?����X�?             @C      D                    �@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @G      H      
             @j#;��h�?*            �P@������������������������       �                     *@I      ^      	            ��@�QA�!�?$             K@J      U                   �?>@�?��?            �E@K      L                ����?�G�z��?             4@������������������������       �                     @M      T      
            �2@     ��?             0@N      O                   "�@�q�q�?	             (@������������������������       �                     @P      Q                   @      �?              @������������������������       �                     @R      S                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @V      W                   F@t���?             7@������������������������       �                     &@X      [                ����?�q�q�?             (@Y      Z                   �?      �?             @������������������������       �                     �?������������������������       �                     @\      ]                   @      �?              @������������������������       �                     �?������������������������       �                     @_      `                   f�@�C��2(�?             &@������������������������       �                     @a      b      	            V�@r�q��?             @������������������������       �                     @������������������������       �                     �?d      m                  @O@`��F:u�?7            �U@e      l                   ��@�Ń��̧?5             U@f      k                   �?r�q��?             (@g      j      
             #@�q�q�?             @h      i                   .@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@������������������������       �        .             R@n      o      
             0@�q�q�?             @������������������������       �                      @������������������������       �                     �?q      L                   6�@P�T���?�           p�@r      �      	            @I�l�~c�?q           �@s      x                   ғ@�����?y            �h@t      u      	            �@ ������?N            �_@������������������������       �        J            �]@v      w                   ��@      �?              @������������������������       �                     @������������������������       �                      @y      z                   �@x�� ���?+            @R@������������������������       �                     @{      �                ���@z�G�z�?)            �Q@|      �                   .@���c���?             J@}      �                   �?t��ճC�?             F@~                         ��@"pc�
�?             &@������������������������       �                     "@������������������������       �                      @�      �                   �?Pa�	�?            �@@������������������������       �        
             3@�      �                   2@@4և���?             ,@�      �                   @z�G�z�?             @������������������������       �                     @�      �      
             '@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     "@�      �                   @      �?              @������������������������       �                     @������������������������       �                     @�      �                   @b�2�tk�?
             2@�      �                   �?      �?             ,@������������������������       �                     @�      �                   @�z�G��?             $@�      �                   �?���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @�      �                   ��@��O,���?�            `y@�      �                   �@��� ?�?i            �f@�      �                  �8@�L:�d�?            �@@�      �                   d�@     ��?	             0@�      �      	            -�@      �?             (@������������������������       �                     "@������������������������       �                     @������������������������       �                     @�      �                   �?.k��\�?             1@�      �                   #@�Q����?             @������������������������       �                     @�      �      	            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     (@�      �                   '@Z���Q��?T            �b@�      �      	            �@�tD�,Y�?O             a@�      �      	            ��@�eP*L��?             F@�      �      
             3@f���M�?             ?@�      �                  @F@8^s]e�?             =@�      �      
             @z�G�z�?             9@�      �                   %@      �?             @������������������������       �                     �?�      �                   ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   @؇���X�?             5@�      �                   $�@      �?              @�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     *@������������������������       �                     @������������������������       �                      @������������������������       �                     *@�      �      	            �@l���?4            @W@�      �                  �K@     ��?#             P@�      �                ����?�NW���?            �J@�      �                   @      �?              @������������������������       �                     @�      �                   %@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                   .@����?�?            �F@�      �                   �?؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     C@�      �                   ԃ@���!pc�?             &@������������������������       �                     @������������������������       �                      @�      �                   �?>���Rp�?             =@�      �                   �@b�2�tk�?             2@�      �                   �?r�q��?             (@������������������������       �                     �?�      �                   �?"pc�
�?             &@������������������������       �                     �?�      �                pff�?ףp=
�?             $@������������������������       �                     "@������������������������       �                     �?�      �                   @r�q��?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     &@�      �                  @@@VUUUUU�?             (@�      �                   �?z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @�      �      
             #@�S�r
>�?�             l@�      �                   0@��o�u<�?5            �T@�      �      	            o�@�;&	���?-            @P@�      �                   @<ݚ)�?             B@�      �                   |�@V�a�� �?             =@�      �                   �?      �?             @������������������������       �                      @�      �                `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?H%u��?             9@������������������������       �                     �?�      �                   @�8��8��?             8@������������������������       �                     (@�      �                   %@r�q��?	             (@�      �                   @�C��2(�?             &@������������������������       �                     @�      �                   �?z�G�z�?             @�      �      
             @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �      
             @����X�?             @������������������������       �                     @�      �      	            ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     =@�      �                   *@�t����?             1@�      �                `ff�?      �?             0@�      �      
             @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     *@������������������������       �                     �?       5      
            �0@�M�Q��?Z            �a@      0                  �2@*a����?>            �X@            	            ��@j���f�?9            �V@                         @�(��w�?            �E@                         l�@և���X�?             @������������������������       �                     @������������������������       �                     @                        �8@O��E�?             B@                         @     ��?
             0@	      
      	            �@�q�q�?             @������������������������       �                      @������������������������       �                     @                         �?ףp=
�?             $@                         2�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @            	            l�@P���Q�?
             4@                         �?      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     0@      %                   @!d���e�?!            �G@      $      	            ��@̂U��?             ?@                         ��@�q�q�?             8@������������������������       �                     �?                         �?�LQ�1	�?             7@                         7@      �?             @������������������������       �                      @������������������������       �                      @                         ĕ@�}�+r��?             3@������������������������       �                     (@       #                ����?؇���X�?             @!      "                ����?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @&      /      
             .@      �?             0@'      (                   .@����X�?
             ,@������������������������       �                     @)      *      
             %@      �?              @������������������������       �                      @+      ,                  �0@�q�q�?             @������������������������       �                     �?-      .                  @B@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @1      2                   @�<ݚ�?             "@������������������������       �                     �?3      4      	            w�@      �?              @������������������������       �                     @������������������������       �                     �?6      E                   @B;��ź�?            �E@7      :                   ��@G���ջ�?             :@8      9                   8�@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@;      >                   `�@     @�?
             0@<      =                    @      �?             @������������������������       �                      @������������������������       �                      @?      @                `ff@VUUUUU�?             (@������������������������       �                     @A      B                    @z�G�z�?             @������������������������       �                     �?C      D      	            �@      �?             @������������������������       �                     @������������������������       �                     �?F      G                   .@������?             1@������������������������       �                      @H      I                  �E@�r����?	             .@������������������������       �                     (@J      K                  �I@�q�q�?             @������������������������       �                      @������������������������       �                     �?M      P                   ��@d(Q���?s             f@N      O      	            ��@d}h���?             ,@������������������������       �                     &@������������������������       �                     @Q      T                   @�G��c�?m            `d@R      S      
            �3@      �?              @������������������������       �                     @������������������������       �                     �?U      ~      	            ��@��<�^�?h            `c@V      g                   �?������?2            �R@W      \      	            ȉ@��s��t�?            �D@X      [      
             @@4և���?
             ,@Y      Z                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@]      ^                   �?������?             ;@������������������������       �                     (@_      d                ����?��S���?
             .@`      c                   @؇���X�?             @a      b                `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @e      f      
            �0@      �?              @������������������������       �                     @������������������������       �                     �?h      s                   l�@߄*�u�?             A@i      j      	            ��@�GN��?             6@������������������������       �                     @k      r                   �?0�����?             2@l      q                   %@�������?             (@m      n                   �?�C��2(�?             &@������������������������       �                     @o      p      
             .@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @t      }                  @J@9��8���?             (@u      |                ���@      �?              @v      w      	            ��@�Q����?             @������������������������       �                     �?x      {                   -@      �?             @y      z                033@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @      �                `ff @��Q�^�?6             T@�      �      	            ��@     ��?*             P@�      �                   �@��k=.��?            �G@�      �                   @և���X�?             @������������������������       �                     @������������������������       �                     @�      �                   !@R���Q�?             D@�      �                033�?`Jj��?             ?@�      �      	            ��@؇���X�?             ,@������������������������       �                     (@������������������������       �                      @������������������������       �                     1@�      �                `ff�?X�<ݚ�?             "@������������������������       �                     @�      �                   �@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     1@�      �      	            �@     ��?             0@�      �                  �A@�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                   ��@$�q-�?	             *@�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     &@�t�bh�h(h+K ��h-��R�(KM�KK��hb�B S       �z@     @y@     �y@     Pv@     �h@      h@      l@     �i@     �h@     �d@      ?@              N@     �A@       @              "@                             �I@     �A@       @             �G@      @                      A@      �?                      @      �?                      @                                      �?                      ;@                              *@      @                      (@                              �?      @                              @                      �?                              @      ?@       @              @      "@      @                               @              @      "@      @              @      @      @               @      @       @               @      @                              @                       @       @                       @                                       @                                       @              �?      �?       @              �?      �?                      �?                                      �?                                       @                      @                      �?      6@       @                      �?      �?                              �?                      �?                      �?      5@      �?              �?                                      5@      �?                      &@      �?                      @                              @      �?                              �?                      @                              $@                      a@     �`@      7@             �V@      ?@       @              ;@      @                      ;@      @                      ;@                                      @                              �?                     �O@      9@       @              C@      4@       @              9@      @       @              (@      @       @                      @                      (@      �?       @               @      �?       @               @      �?                              �?                       @                                               @              $@                              *@                              *@      .@                      @      &@                      @      $@                      @       @                      �?       @                               @                      �?                               @                                       @                       @      �?                              �?                       @                               @      @                               @                       @       @                       @                                       @                      9@      @                      .@      @                      @      @                      @                               @      @                              @                       @      �?                              �?                       @                              $@      �?                      $@                                      �?                      $@                             �G@     @Y@      5@              =@     �U@      &@              *@      @@      @              (@      7@      @               @      6@      @               @       @      �?               @      @      �?              @              �?                              �?              @                              @      @                      @                                      @                              @                              ,@      @                              �?                      ,@       @                      $@                              @       @                      @                                       @              @      �?      @               @                               @      �?      @               @      �?                              �?                       @                                              @              �?      "@                      �?      @                              @                      �?                                      @                      0@      K@      @              .@      @                      @                              "@      @                      �?      @                              @                      �?                               @                              �?     �I@      @              �?     �@@                              ?@                      �?       @                      �?                                       @                              2@      @                      @       @                      @      �?                       @                               @      �?                              �?                       @                                      �?                      ,@       @                      @       @                      @      �?                              �?                      @                                      �?                      @                      2@      .@      $@              1@                              �?      .@      $@              �?      &@      �?              �?      �?                              �?                      �?                                      $@      �?                              �?                      $@                              @      "@                      @      "@                               @                      @      �?                      �?                               @      �?                       @                                      �?                      �?                              :@      h@     �i@              (@     �W@     �S@              @      B@      @              @       @                      �?                               @       @                       @                                       @                      �?      A@      @              �?      9@      @                      0@       @                      (@                              @       @                               @                      @                      �?      "@      @              �?                                      "@      @                       @                              �?      @                              @                      �?      �?                              �?                      �?                              "@                       @     �M@      R@              �?      =@      4@              �?      .@      @              �?      "@      @              �?       @      @              �?              @                              @              �?                                       @                              @                              @       @                       @      �?                       @                                      �?                      @      �?                      @                                      �?                      ,@      ,@                      &@      @                      @      @                      �?      @                      �?                                      @                      @      �?                      @                                      �?                      @                              @       @                      @       @                       @                              �?       @                      �?                                       @                              @              @      >@      J@               @      @      9@               @      @      8@                              "@               @      @      .@               @       @                               @                       @                                      �?      .@                              (@                      �?      @                      �?                                      @                      @      �?                      �?      �?                      �?                                      �?                       @                      @      8@      ;@              @      8@      1@               @      "@      *@                              �?               @      "@      (@               @       @       @                               @               @       @                       @       @                               @                       @                                      @                              �?      $@                              @                      �?      @                      �?                                      @              @      .@      @                       @                      @      @      @              @      �?      @                              @              @      �?      �?              @              �?              @                                              �?                      �?                              @                                      $@              ,@     �X@     @_@              ,@     �W@      E@                      ;@      @                      5@      �?                      5@                                      �?                      @      @                      @       @                      @                               @       @                               @                       @                                       @              ,@     �P@     �B@              *@      B@       @               @      >@       @               @      @                       @                                      @                              :@       @                      *@       @                      "@                              @       @                      @      �?                      @                                      �?                      �?      �?                      �?                                      �?                      *@                      &@      @                      @                              @      @                              @                      @      @                              �?                      @       @                       @       @                       @                                       @                      @                              �?      ?@     �A@                              *@              �?      ?@      6@              �?      >@      (@                      &@      "@                      @                              @      "@                      @      @                              @                      @      �?                      @                               @      �?                              �?                       @                                      @              �?      3@      @                      &@                      �?       @      @                      �?      @                      �?                                      @              �?      @                      �?                                      @                              �?      $@                              @                      �?      @                              @                      �?                              @     �T@                       @     �T@                       @      $@                       @      �?                      �?      �?                      �?                                      �?                      �?                                      "@                              R@                       @      �?                       @                                      �?     @m@     `j@      g@      c@     �j@     �d@     @^@     @Z@     �f@      3@                      _@       @                     �]@                              @       @                      @                                       @                      L@      1@                              @                      L@      ,@                     �F@      @                     �D@      @                      "@       @                      "@                                       @                      @@      �?                      3@                              *@      �?                      @      �?                      @                              �?      �?                              �?                      �?                              "@                              @      @                              @                      @                              &@      @                      @      @                      @                              @      @                      @       @                               @                      @                                      @                      @                              @@     �b@     @^@     @Z@      =@     �L@      P@      @@      "@      1@      @      @      "@      @      @              "@              @              "@                                              @                      @                              *@      �?      @              �?      �?      @                              @              �?      �?                      �?                                      �?                      (@                      4@      D@      N@      =@      4@      B@     �M@      6@      4@      8@                      4@      &@                      4@      "@                      4@      @                       @       @                      �?                              �?       @                               @                      �?                              2@      @                      @      @                      �?      @                      �?                                      @                      @                              *@                                      @                               @                              *@                              (@     �M@      6@              (@      J@                      @     �H@                      @      @                              @                      @       @                      @                                       @                      �?      F@                      �?      @                      �?                                      @                              C@                       @      @                              @                       @                                      @      6@                      @      &@                       @      $@                              �?                       @      "@                      �?                              �?      "@                              "@                      �?                              @      �?                              �?                      @                                      &@              @      �?      @              @      �?                      @                                      �?                                      @      @     �V@     �L@     @R@              D@      &@      ?@              9@      &@      =@              9@      &@                      7@      @                      �?      @                               @                      �?      �?                              �?                      �?                              6@      @                              �?                      6@       @                      (@                              $@       @                      $@      �?                      @                              @      �?                       @      �?                       @                                      �?                       @                                      �?                       @      @                              @                       @      �?                       @                                      �?                                      =@              .@               @              .@              �?               @              �?               @                                              �?              *@                                              �?      @     �I@      G@      E@      �?      A@      E@      6@      �?      A@     �A@      4@      �?     �@@      "@                      @      @                      @                                      @              �?      >@      @                      &@      @                       @      @                       @                                      @                      "@      �?                       @      �?                              �?                       @                              @                      �?      3@                      �?      @                      �?                                      @                              0@                              �?      :@      4@              �?      4@      $@              �?      4@      @              �?                                      4@      @                       @       @                       @                                       @                      2@      �?                      (@                              @      �?                      �?      �?                      �?                                      �?                      @                                      @                      @      $@                      @      $@                              @                      @      @                       @                               @      @                              �?                       @      @                              @                       @                               @                              @       @                              �?                      @      �?                      @                                      �?       @      1@      @      4@       @      *@      @      @              "@      �?                              �?                      "@                       @      @      @      @       @               @               @                                               @                      @      �?      @                              @              @      �?                      �?                              @      �?                      @                                      �?                      @              *@               @                               @              *@                              (@               @              �?               @                                              �?      6@      F@     �O@      H@                      &@      @                      &@                                      @      6@      F@      J@     �F@              �?              @                              @              �?                      6@     �E@      J@      C@      6@      E@      &@              *@      5@      @              *@      �?                       @      �?                              �?                       @                              &@                                      4@      @                      (@                               @      @                      �?      @                      �?      �?                              �?                      �?                                      @                      @      �?                      @                                      �?              "@      5@      @              @      0@      �?              @                              �?      0@      �?              �?      $@      �?                      $@      �?                      @                              @      �?                      @                                      �?              �?                                      @                      @      @      @              @      �?      @              �?      �?      @              �?                                      �?      @                      �?      �?                              �?                      �?                                       @              @                                      @                              �?     �D@      C@                      C@      :@                      C@      "@                      @      @                      @                                      @                      A@      @                      =@       @                      (@       @                      (@                                       @                      1@                              @      @                              @                      @      �?                      @                                      �?                              1@              �?      @      (@              �?       @                               @                      �?                                      �?      (@                      �?      �?                              �?                      �?                                      &@�t�bub�H6     hhubh)��}�(hhhhhNhKhKhG        hh$hNhJ�v}hG        hNhG        hHKhIKhJh(h+K ��h-��R�(KK��hb�C               �?       @      @�t�bhVhghQC       ���R�hkKhlhoKh(h+K ��h-��R�(KK��hQ�C       �t�bK��R�}�(hKhyM�hzh(h+K ��h-��R�(KM���h��B��         �                   �?��6���?�            �@       i                   !@���r`��?           P�@       $                   @+��K���?�           ��@       �                 ���@dF���?J           p�@       �                    %@�8-s��?           pz@       	                    @R�n���?�             r@                           ��@�q�q�?             "@������������������������       �                     @������������������������       �                     @
       k                    Ė@�2�8���?�            pq@       0                    �?@���d�?p            `f@       #                    �?��:��?1            @U@                           #@
dq"��?%            �O@������������������������       �                     @       "       
            �3@8>�ݜ��?"            �M@       !                    @j�V��?!            �L@                           d�@�!���O�?             �K@              	            �@և���X�?             @������������������������       �                     @������������������������       �                     @              	            ^�@VUUUU��?             H@������������������������       �                    �B@                           �?�C��2(�?
             &@������������������������       �                      @                           �@h/�����?	             "@������������������������       �                     @                           @O@      �?             @                           @z�G�z�?             @                          @H@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                      @$       +                   �;@J���#�?             6@%       &       
             @      �?              @������������������������       �                      @'       *                    @      �?             @(       )       
            �0@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @,       -       	            ��@T�r
^N�?             ,@������������������������       �                      @.       /       
             +@r�q��?             @������������������������       �                     @������������������������       �                     �?1       f                    >�@i��a��??            �W@2       e                    ,�@Y\���?:            �U@3       R                   @G@<rN?��?9            �T@4       G                    p�@�h$��W�?&             N@5       6       	            <�@�Y����?             E@������������������������       �                     (@7       @                    �?���� C�?             >@8       =       	            a�@@�0�!��?
             1@9       :                    @"pc�
�?             &@������������������������       �                     @;       <                    @      �?             @������������������������       �                      @������������������������       �                      @>       ?       	            ��@�q�q�?             @������������������������       �                     @������������������������       �                      @A       F       	            6�@�	j*D�?             *@B       E                    .@z�G�z�?             @C       D       
             )@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @H       I                    @x�5?,�?             2@������������������������       �                     �?J       M       	            F�@:���I�?             1@K       L                    @���Q��?             @������������������������       �                      @������������������������       �                     @N       Q                   �6@�8��8��?             (@O       P                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@S       \                 pff�?X��t��?             7@T       W                    �?      �?              @U       V       
             *@      �?             @������������������������       �                     @������������������������       �                     �?X       [                    ��@      �?             @Y       Z                 ����?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?]       d                    @N贁N�?             .@^       a                   �M@�m۶m��?             ,@_       `                    @�8��8��?	             (@������������������������       �                     &@������������������������       �                     �?b       c       
             @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     @g       h       	             �@      �?              @������������������������       �                     �?i       j                    �?؇���X�?             @������������������������       �                     �?������������������������       �                     @l       �                   @F@����x��?D             Y@m       n                    `�@���~�?6            �R@������������������������       �                     @o       �                    @�[��_�?4            �Q@p              	            �@����N�?"            �H@q       v                    �?�&���?             >@r       u       
             #@j�V���?             &@s       t                    (@�����H�?             "@������������������������       �                     �?������������������������       �                      @������������������������       �                      @w       z                    �?�����?             3@x       y       	            �@      �?             @������������������������       �                     @������������������������       �                     @{       |       
             +@�θ�?             *@������������������������       �                     @}       ~                    <@      �?             @������������������������       �                     @������������������������       �                     @�       �                    �?D�n�3�?             3@�       �                    �?���Q��?             $@�       �       
             *@����X�?             @������������������������       �                      @������������������������       �                     @�       �       	            c�@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	            &�@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    x�@��!pc�?             6@�       �                    �?      �?              @�       �                    �?      �?             @������������������������       �                      @�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?�       �                     @      �?             @������������������������       �                     �?������������������������       �                     @�       �                    �?X�Cc�?             ,@�       �                    ��@      �?             $@�       �       	            ��@      �?              @������������������������       �                     @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �                   �N@�������?             9@�       �       	            ��@t���?             7@�       �                    �@�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    �?P���Q�?             4@�       �                   �L@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �        	             1@������������������������       �                      @�       �                   �M@�w7lh�?O            �`@�       �       
             @`�BE��?I             _@�       �                 033�?����X�?             @�       �       	            �@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�       �                    �?UQ[Z��?E            @]@�       �       	            ��@S�K�0��?            �E@�       �                    ��@     ��?             0@�       �                    @      �?              @������������������������       �                     @�       �                    �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                 033�?�����H�?             ;@�       �       	            ��@�z�G��?             $@�       �                    4@���Q��?             @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �        
             1@�       �                    �?\� sAr�?)            �R@�       �                    �?Z;����?             A@�       �                   �K@�n���?             "@�       �                    �?�8��8��?             @������������������������       �                     @�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�       �                    �?jM��?             9@�       �                    �?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �                    @��|���?             6@������������������������       �                     @�       �       	            `�@�W�3��?             3@�       �                    v�@�����H�?             "@������������������������       �                      @������������������������       �                     �?�       �                    0@��(\���?             $@�       �       	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                 ���@      �?              @������������������������       �                     @������������������������       �                     �?�       �                    @{�G�z�?             D@�       �       	            �@�ӭ�a��?             2@�       �                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     .@�       �       	            ��@�GN��?             6@�       �                    )@�IєX�?	             1@�       �                    J@      �?             @�       �                    :@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                     @�       �       	            |�@���k���?             &@������������������������       �                      @�       �       
             /@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �       	             �@���B[��?C            �Y@�       �                    %@��V�I��?             �G@�       �       	            f�@�5��?             ;@������������������������       �                     @�       �                    @z�G�z�?             4@�       �                    �?�����H�?             2@�       �                    l�@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     (@������������������������       �                      @�       �       	            ��@      �?             4@������������������������       �                     &@�       �                    H�@X�<ݚ�?             "@�       �       
             $@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�                          @�X�C�?#             L@�                          @
ףp=
�?             4@                          �?      �?             @                      033@VUUUUU�?             @������������������������       �                     �?            	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @                        �8@/����?             ,@      	                   @      �?             @������������������������       �                     �?
                         1@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@                      ���@�q�q�?             B@            	            ��@�q�q�?             8@                         �?ףp=
�?             4@������������������������       �                     �?                        �6@�}�+r��?
             3@                         ��@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@            
             '@      �?             @������������������������       �                     @������������������������       �                     �?                          @��8��8�?             (@                        �0@�Q����?             @������������������������       �                     @            
             ,@      �?              @������������������������       �                     �?������������������������       �                     �?       !                    �@����X�?             @������������������������       �                     �?"      #                   /@r�q��?             @������������������������       �                     @������������������������       �                     �?%      &                   t�@�����L�?`            �a@������������������������       �                     @'      B      	            �@�Qߛ�F�?^             a@(      ;                   #@؇���X�?&             L@)      .                   �?��Q��?             4@*      -      
             &@�q�q�?             @+      ,                `ff�?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?/      4                   �?�t����?             1@0      3      
             -@�q�q�?             @1      2                   �?z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?5      :                   @�C��2(�?             &@6      7                   �?      �?             @������������������������       �                      @8      9                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @<      A                   �?������?             B@=      >                   �?r�q��?             @������������������������       �                     @?      @                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     >@C      Z                   �?`��`s�?8            @T@D      Y      	            Щ@�8��8��?!             H@E      L                   ?@(N:!���?            �A@F      I                   �?�r����?             .@G      H                   �?�C��2(�?             &@������������������������       �                     $@������������������������       �                     �?J      K                   ��@      �?             @������������������������       �                     �?������������������������       �                     @M      T                  @D@��Q��?             4@N      S                  �A@����X�?             @O      P      
             @�q�q�?             @������������������������       �                     �?Q      R                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @U      X                   2@8�Z$���?	             *@V      W      	            ��@�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?������������������������       �                     *@[      d      	            �@cڟXǰ�?            �@@\      c                033@�8��8��?
             (@]      b      	            �@      �?              @^      _      	            ��@�q�q�?             @������������������������       �                     @`      a                   @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @e      h      
             @�����?             5@f      g                   @�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �        	             .@j      �                   �@*!c`vu�?^            �a@k      n                   �?�:���?            �G@l      m      
            �1@���Q��?             @������������������������       �                     @������������������������       �                      @o      r                   D�@��{�~�?             E@p      q                033@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @s      z      	            *�@���{���?            �@@t      y                   �?��S�ۿ?	             .@u      x                  @N@      �?             @v      w      	            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     &@{      �      
            �2@VUUUUU�?             2@|      �      	            �@VUUUUU�?             .@}      �                   �?      �?              @~                         @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @�      �                  @@@և���X�?             @������������������������       �                     @�      �      	            >�@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �      	            �@O��1��?@            �W@�      �      	            ��@61��?0            �Q@�      �                   �?1X�ܐ^�?#            �G@�      �                `ff�?�X�<ݺ?             2@������������������������       �                     ,@�      �                   ��@      �?             @������������������������       �                     @������������������������       �                     �?�      �                   .@CbΊx�?             =@�      �                   '@      �?              @�      �                   @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                   ��@d��b��?             5@������������������������       �                     @�      �                   +@     @�?             0@�      �                   @      �?              @������������������������       �                     �?�      �                   '@0�����?             @�      �      
             @      �?             @������������������������       �                      @�      �      	            H�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                  @H@      �?              @������������������������       �                     @�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   /@�nkK�?             7@������������������������       �        
             3@�      �                   @      �?             @������������������������       �                      @�      �                   ��@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   *�@`2U0*��?             9@�      �                   @؇���X�?             @�      �                   #@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     2@�      L                   @m�~��?�           ��@�                         @��{ri`�?�            �o@�      �                  @B@;�yz7�?S            �`@�      �                   @�G�zT�?0             T@�      �                   �?     x�?*             P@�      �                   �?cڟXǰ�?            �@@�      �                   �@Ra���i�?             6@�      �                   �?�ӭ�a��?
             2@�      �                   �?�$I�$I�?             @�      �                   @      �?             @������������������������       �                     �?�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     &@�      �                  �2@      �?             @������������������������       �                      @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   @"pc�
�?             &@�      �                  �A@X�<ݚ�?             "@�      �                   `�@؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                      @�      �      	            ؈@�-��?             ?@������������������������       �                     &@�      �                   �?�(\����?             4@�      �      	            Ӣ@�8��8��?             @������������������������       �                      @�      �                   Ƒ@      �?             @������������������������       �                     �?������������������������       �                     @�      �                ����?������?             ,@������������������������       �                      @�      �      
             #@      �?
             (@�      �                   @{�G�z�?             @�      �                  �8@�q�q�?             @������������������������       �                     �?�      �      
             @      �?              @������������������������       �                     �?������������������������       �                     �?�      �      	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   @؇���X�?             @������������������������       �                     @������������������������       �                     �?�      �                   2@     ��?             0@�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @�      �                   �?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@�                         �?ƵHPS!�?#             J@�      �                   J@:J�����?             :@�      �                @33�?|�l�]�?             1@������������������������       �                      @�      �                   G@$߼�x�?             .@�      �                   �?      �?              @������������������������       �                     @�      �                   �?      �?             @������������������������       �                      @�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   D�@և���X�?             @�      �      	            ��@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                      @                          �?X�<ݚ�?             "@������������������������       �                     @            
             @{�G�z�?             @������������������������       �                      @                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @      
                  �F@���3�E�?             :@      	                   ��@ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@                         0�@      �?             0@            	            �@؇���X�?             @������������������������       �                     @������������������������       �                     �?                         M@�q�q�?             "@            	            צ@���Q��?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @            	            ̖@�vCu��?K            �^@                         t�@�?�'�@�?             C@            	            x�@�IєX�?             A@������������������������       �                     ;@                         @����X�?             @������������������������       �                     @������������������������       �                      @                         �?      �?             @������������������������       �                     �?������������������������       �                     @      =                  �H@��t�_�?1            @U@      2      	            A�@��IB���?%            @P@       !                   !@�^�����?            �C@������������������������       �                     @"      1      
            �1@���Er�?             A@#      0                   @w���<�?             ?@$      +                `ff @�8��8��?             8@%      *      	            �@B{	�%��?	             2@&      )                   H�@      �?             0@'      (                   (�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �                      @,      /                   @r�q��?             @-      .      	            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @������������������������       �                     @3      4                   �?�	j*D�?             :@������������������������       �                     $@5      8                   �?      �?             0@6      7                  @E@z�G�z�?             @������������������������       �                     @������������������������       �                     �?9      <                   @���|���?             &@:      ;                  �0@և���X�?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @>      E      
             '@��(\���?             4@?      @      
             @{�G�z�?             $@������������������������       �                     @A      D      	            �@�$I�$I�?             @B      C                  �J@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @F      G                   �?��(\���?             $@������������������������       �                     @H      I                   �?      �?             @������������������������       �                      @J      K                   @      �?              @������������������������       �                     �?������������������������       �                     �?M      ~                  �0@���J��?F           ��@N      W                   @�I �\��?@           h�@O      �                  �=@�0��7��?           �{@P      �                   �?��F���?�             j@Q      �                  �1@�gZ���?8            �S@R      �      
            �0@'&��|��?/            �P@S      h                   �?�e�c]��?%             I@T      U                   �?
ц�s�?             :@������������������������       �                     @V      [                   4�@"pc�
�?             6@W      X                   �?z�G�z�?             @������������������������       �                     @Y      Z                   .@      �?              @������������������������       �                     �?������������������������       �                     �?\      ]                   �?ҳ�wY;�?             1@������������������������       �                      @^      e                   �?��S���?	             .@_      b                   @�q�q�?             (@`      a      	            ؔ@؇���X�?             @������������������������       �                     �?������������������������       �                     @c      d                  �6@���Q��?             @������������������������       �                     @������������������������       �                      @f      g      	            ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @i      v                   �?      �?             8@j      s                   -@�g���e�?             &@k      r                   �?      �?              @l      q                   @      �?             @m      n      
             *@z�G�z�?             @������������������������       �                      @o      p                   d�@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @t      u      	            ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @w      �      	            ŧ@�1G����?             *@x      }                ����?��E���?             "@y      |                   �?      �?             @z      {      
             @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     �?~            	            *�@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �      	            Κ@k��\��?
             1@������������������������       �                     "@�      �                   �?      �?              @�      �                   �?{�G�z�?             @�      �                   ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   @VUUUUU�?	             (@�      �                   �?      �?             @������������������������       �                     �?������������������������       �                     @�      �      	            @      �?              @�      �                   �?؇���X�?             @�      �                   �?r�q��?             @������������������������       �                     �?�      �                  �4@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?�      �                   /@,�wɃ�?P            @`@�      �                   -@ܝ��.4�?O            @_@�      �                   )@��#�]�?7            �V@�      �                   <�@��ǒ��?(             O@�      �                `ff�?�$�_�?
             3@������������������������       �                     @�      �                   �?     @�?	             0@������������������������       �                     @�      �      	            ��@��8��8�?             (@������������������������       �                     @�      �                   2@r�q��?             @������������������������       �                     @������������������������       �                     �?�      �                   \�@ޓtf���?            �E@�      �                033�?�����H�?             "@������������������������       �                     @�      �      
              @      �?              @������������������������       �                     �?������������������������       �                     �?�      �      
             @�������?             A@�      �                   �?r�q��?             @�      �      	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �      
             %@����S��?             <@�      �                   �?r�q��?             @������������������������       �                     @�      �                   #@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   �?}��7�?             6@�      �                   @b���i��?	             &@�      �                   @      �?              @������������������������       �                     �?������������������������       �                     �?�      �      	            ܔ@�n���?             "@������������������������       �                     @�      �      	            ��@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                pff�?�g���e�?             &@������������������������       �                     @�      �                   ��@�8��8��?             @�      �                    @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                  �5@�����\�?             =@�      �                   �?���QI�?             9@�      �      	            �@�8��8��?             (@������������������������       �                     "@�      �                   @�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �                   �?&�q-�?             *@�      �      	            �@؇���X�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �                   �?�������?             A@�      �      	            ϡ@�eP*L��?             &@������������������������       �                     @������������������������       �                     @�      �                   p�@�[")�i�?             7@�      �      	            Z�@�'}�'}�?             .@�      �                   !@ףp=
�?             $@������������������������       �                      @�      �                   
�@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                  �0@���Q��?             @������������������������       �                     @������������������������       �                      @�      �                   @      �?              @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @�      �      
             @=��h[�?�             m@�      �      	            H�@     ��?
             0@�      �                   �?���|���?             &@������������������������       �                     �?�      �                   �?�z�G��?             $@������������������������       �                     @�      �                   �?      �?             @������������������������       �                     @������������������������       �                     @������������������������       �                     @�      P      	            z�@61j�)�?             k@�      C                   ��@7w,k�.�?`            `c@�      .                  �0@���y&�?Q            @`@�                         �?/�w�$�?=            �X@�      
      
            �2@��!pc�?            �@@�                         А@x9/���?             <@�      �                ����?     @�?             0@������������������������       �                     @�                         �G@      �?             (@�      �                   ��@և���X�?             @������������������������       �                     @������������������������       �                     @                        �K@���Q��?             @������������������������       �                     @������������������������       �                      @                         �?r�q��?             (@������������������������       �                     �?      	                   �?�C��2(�?             &@                         !@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @            	            �@z�G�z�?             @������������������������       �                     �?������������������������       �                     @      -                   @R/s?o�?$            @P@                         �?���)�?!            �M@                         ��@�������?             (@                         @�C��2(�?             &@                         ��@r�q��?             @������������������������       �                     @                         �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     �?                          �?��[�p�?            �G@            
             1@     ��?             0@                      pff@.y0��k�?             *@                         .@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?������������������������       �                     �?������������������������       �                     @!      ,                033�?�[���q�?             ?@"      %      	            �@"��u���?             9@#      $                   �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@&      '                   l�@�r����?             .@������������������������       �                     (@(      )                   �?�q�q�?             @������������������������       �                     �?*      +                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                     @/      8      
             -@     ��?             @@0      1                   �?����X�?             5@������������������������       �                      @2      3                   �?���y4F�?             3@������������������������       �                      @4      5                   �?�t����?	             1@������������������������       �                     "@6      7                   H@      �?              @������������������������       �                      @������������������������       �                     @9      <      
             /@}��7�?             &@:      ;                  �G@      �?             @������������������������       �                      @������������������������       �                      @=      B      	            �@�$I�$I�?             @>      ?      
            �1@�q�q�?             @������������������������       �                     �?@      A                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @D      I                   X�@��A�f�?             9@E      H      	            0�@޾�z�<�?             *@F      G                  �2@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     $@J      M                033�?      �?             (@K      L                   @z�G�z�?             @������������������������       �                     @������������������������       �                     �?N      O      	            ��@؇���X�?             @������������������������       �                     �?������������������������       �                     @Q      V                   @�@`Jj��?             O@R      S                   (@\-��p�?             =@������������������������       �                     ,@T      U                   "@������?             .@������������������������       �                     &@������������������������       �                     @������������������������       �                    �@@X      [      	            h�@*�jE���?/            �T@Y      Z                   �?�#-���?            �A@������������������������       �                     @������������������������       �                     @@\      m                ����?�q�q��?              H@]      f                   �?�<ݚ�?             2@^      _      
             @      �?              @������������������������       �                     �?`      e                   P�@�$I�$I�?             @a      b                   �?      �?             @������������������������       �                     �?c      d                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @g      l                   @�z�G��?             $@h      k                `ff�?���Q��?             @i      j                   0@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @������������������������       �                     @n      u                   �?�8��8��?             >@o      p      	             �@�$I�$I�?             @������������������������       �                     @q      t                   �?�q�q�?             @r      s                   |�@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?v      w                033�?\1�K36�?             7@������������������������       �                     "@x      }      	            �@T�r
^N�?             ,@y      z                   �?r�q��?             @������������������������       �                     @{      |      
            �0@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @      �                   @��(\���?             $@������������������������       �                     �?�      �      
             #@�����H�?             "@������������������������       �                     �?������������������������       �                      @�t�bh�h(h+K ��h-��R�(KM�KK��hb�B`p        y@      y@     Py@     �x@     �g@      g@     �k@     �j@     �d@     @a@     `f@      g@     �]@     �]@     �a@     �b@      W@     �V@      \@      `@     @T@     �L@     �R@      S@      @      @                              @                      @                             �R@      K@     �R@      S@     �O@      >@      H@      C@      D@      .@      3@      &@     �B@      @      *@      @                      @             �B@      @      "@      @     �B@      @      "@      @     �B@      @      @      @              @      @                      @                                      @             �B@      @      @      @     �B@                                      @      @      @               @                              �?      @      @                              @              �?      @      �?              �?      @                      �?       @                      �?                                       @                               @                                      �?                       @                                       @      @       @      @      @      @              �?      @       @                              �?              �?      @      �?              �?              �?                                              �?                                      @               @      @      �?               @                                      @      �?                      @                                      �?      7@      .@      =@      ;@      6@      .@      7@      :@      3@      .@      7@      :@      .@      (@      &@      6@      (@      "@      $@      &@      (@                                      "@      $@      &@              "@      @       @              "@       @                      @                               @       @                       @                                       @                              @       @                      @                                       @                      @      "@                      @      �?                      �?      �?                              �?                      �?                              @                                       @      @      @      �?      &@              �?                      @       @      �?      &@      @       @                               @                      @                                              �?      &@                      �?       @                               @                      �?                                      "@      @      @      (@      @       @      �?      �?      @                      �?      @                              @                      �?               @      �?              �?       @      �?                              �?                       @                                                      �?       @       @      &@               @      �?      &@              �?              &@                              &@              �?                              �?      �?                              �?                      �?                                      �?                      @                              �?              @      �?      �?                                              @      �?                              �?                      @              (@      8@      :@      C@      &@      6@      7@      3@                              @      &@      6@      7@      .@       @      5@      (@       @       @      5@      �?               @       @      �?                       @      �?                              �?                       @                       @                              @      *@                      @      @                      @                                      @                      @      $@                              @                      @      @                              @                      @                                              &@       @                      @      @                       @      @                       @                                      @                       @      �?                       @                                      �?                      @       @                      @                                       @      @      �?      &@      @      @      �?       @       @              �?       @      �?                       @                      �?              �?              �?                                              �?      @                      �?                              �?      @                                              "@      @                      @      @                      @      @                      @                                      @                       @                              @              �?       @      @      3@      �?              @      3@      �?               @                               @              �?                                              �?      3@                      �?       @                               @                      �?                                      1@               @                      &@     �@@      C@     �J@      "@      ?@      ?@     �J@              @               @               @               @               @                                               @              @                      "@      :@      ?@     �I@      @      "@      @      8@      @      "@                      @      �?                      @                              �?      �?                      �?                                      �?                               @                                      @      8@                      @      @                      @       @                               @                      @                                      @                              1@       @      1@      <@      ;@      �?      0@      $@      @              @       @      @              @       @      �?              @                                       @      �?                              �?                       @                                      @      �?      *@       @      @              �?               @                               @              �?                      �?      (@       @      �?              @                      �?      "@       @      �?      �?       @                               @                      �?                                      �?       @      �?                      �?      �?                      �?                                      �?              �?      @                              @                      �?                      �?      �?      2@      4@      �?               @      .@      �?               @              �?                                               @                                      .@              �?      0@      @              �?      0@                      �?      @                      �?      �?                              �?                      �?                                       @                              *@                                      @       @       @      @               @                                       @      @                              @                       @                      :@      =@      <@      4@      :@      5@                      &@      0@                      @                              @      0@                       @      0@                       @      @                       @                                      @                              (@                       @                              .@      @                      &@                              @      @                      @      �?                              �?                      @                                      @                               @      <@      4@              @      @      &@              @      �?      �?              �?      �?      �?                      �?                      �?              �?              �?                                              �?              @                              �?      @      $@              �?      @                              �?                      �?       @                      �?                                       @                                      $@              @      8@      "@               @      3@      @               @      2@                      �?                              �?      2@                      �?      @                              @                      �?                                      ,@                              �?      @                              @                      �?                      �?      @      @              �?      @      �?                      @                      �?              �?              �?                                              �?                       @      @                      �?                              �?      @                              @                      �?              H@      3@     �C@      B@                      @              H@      3@      A@      B@      H@       @                      *@      @                      �?       @                      �?      �?                              �?                      �?                                      �?                      (@      @                       @      @                      �?      @                      �?                                      @                      �?                              $@      �?                      @      �?                       @                              �?      �?                              �?                      �?                              @                             �A@      �?                      @      �?                      @                               @      �?                       @                                      �?                      >@                                      &@      A@      B@              @      :@      .@              @      :@       @                      *@       @                      $@      �?                      $@                                      �?                      @      �?                              �?                      @                      @      *@                      @       @                      �?       @                              �?                      �?      �?                      �?                                      �?                      @                               @      &@                      �?      &@                      �?                                      &@                      �?                                              *@              @       @      5@              @      @       @              @       @       @              @               @              @                              �?               @              �?                                               @                       @                              @                               @      3@                       @      @                       @                                      @                              .@      8@      G@     �E@      =@      .@      .@      ,@      @               @      @                              @                       @                      .@      *@      &@      @              @      @                      @                                      @              .@       @      @      @      ,@      �?                      @      �?                      �?      �?                              �?                      �?                               @                              &@                              �?      @      @      @      �?      @      @      @      �?      @                      �?       @                      �?                                       @                              @                                      @      @                      @                              �?      @                      �?                                      @                      @              "@      ?@      =@      :@      "@      ?@      <@       @      "@      ?@      @      �?              1@      �?                      ,@                              @      �?                      @                                      �?              "@      ,@      @      �?      @      �?      @                      �?      @                      �?                                      @              @                              @      *@       @      �?              @                      @       @       @      �?      @      �?       @                              �?              @      �?      �?               @      �?      �?               @                                      �?      �?                      �?                                      �?              @                                      @              �?              @                              �?              �?                              �?              �?                                      6@      �?                      3@                              @      �?                       @                              �?      �?                              �?                      �?                              �?      8@                      �?      @                      �?      �?                              �?                      �?                                      @                              2@     �j@      k@     �f@     `f@      T@     �T@     �F@     �G@     �F@     �I@      $@      :@      @@     �A@      @      @      5@      ?@      @      @       @      5@      @              @      .@       @               @      .@      �?               @      @      �?               @      �?      �?                      �?                       @              �?                              �?               @                                      @                              &@                      @              �?               @                              �?              �?                              �?              �?                              @      @       @              �?      @       @              �?      @                      �?                                      @                                       @               @                              *@      $@      @      @      &@                               @      $@      @      @               @      �?      @               @                                      �?      @                      �?                                      @       @       @       @       @                       @               @       @               @       @       @              �?       @      �?                      �?                              �?      �?                              �?                      �?                                      �?              �?              �?                                              �?              @              �?              @                                              �?      &@      @              �?              @              �?                              �?              @                      &@      �?                              �?                      &@                              *@      0@      @      4@      @      (@      @      @      @      @      �?      @               @                      @      @      �?      @       @      @      �?      �?              @                       @              �?      �?       @                                              �?      �?                      �?                                      �?      @                      @      @                       @      @                                                       @                               @      �?      @       @                      @                      �?       @       @                               @              �?       @                      �?                                       @                      @      @              .@      �?                      "@      �?                                                      "@      @      @              @      @      �?                      @                                      �?                              @              @              @               @              @                                               @                              @     �A@      @@     �A@      5@     �@@      @                      @@       @                      ;@                              @       @                      @                                       @                      �?      @                      �?                                      @                       @      ;@     �A@      5@       @      .@      >@      2@       @      .@      6@                      @                       @      $@      6@               @      @      6@               @      @      .@               @       @      ,@               @              ,@               @              �?                              �?               @                                              *@                       @                              @      �?                      �?      �?                      �?                                      �?                      @                                      @                      @                                       @      2@                              $@                       @       @                      @      �?                      @                                      �?                      @      @                      @      @                              @                      @                                      @              (@      @      @              @      @       @              @                              �?      @       @              �?      @                      �?                                      @                                       @               @      �?      �?              @                               @      �?      �?               @                                      �?      �?                              �?                      �?             �`@     �`@     @a@     �`@     ``@     �`@      a@      _@     @X@     @]@     �]@     �[@      P@     �O@     �F@     �B@      9@      .@      7@      0@      2@      &@      6@      0@      "@       @      4@      *@      @              (@       @                              @      @              (@      @      @                      �?      @                              �?                      �?      �?                                                      �?       @              (@      @                       @               @              $@      @      �?               @      @      �?              @              �?                                              @                               @      @                              @                       @              �?               @              �?                                               @              @       @       @      @      �?      @      @              �?      @      �?              �?      @      �?              �?      @                               @                      �?       @                               @                      �?                                              �?                       @                              �?       @                      �?                                       @               @      �?      @      @       @      �?      @      �?       @              �?      �?       @                      �?       @                                                      �?                      �?                      �?      @                      �?                                      @                                      @      "@      @       @      @      "@                                      @       @      @               @       @      �?               @              �?               @                                              �?                       @                      �?               @              �?                                               @      @      @      �?              �?      @                      �?                                      @                      @      �?      �?              @      �?                      @      �?                      �?                              @      �?                      @                                      �?                      �?                                              �?             �C@      H@      6@      5@     �C@     �E@      6@      5@     �B@      <@      ,@      (@      4@      1@      ,@      &@      $@               @      �?                      @              $@              @      �?      @                              @              @      �?      @                                              @      �?                      @                                      �?      $@      1@      @      $@               @      �?                      @                              �?      �?                      �?                                      �?              $@      "@      @      $@      �?      @                      �?      �?                      �?                                      �?                              @                      "@      @      @      $@      @              �?              @                              �?              �?                              �?              �?                              @      @      @      $@      @      �?      @      @              �?              �?                              �?              �?                      @              @       @      @                                              @       @                      @                                       @              @      �?      @                              @              @      �?       @              @      �?                              �?                      @                                               @      1@      &@              �?      1@      @              �?      &@      �?                      "@                               @      �?                              �?                       @                              @      @              �?      @                      �?      @                                                      �?              @                              @                       @      .@       @      "@              @      @                      @                                      @               @      "@      @      "@      �?      "@      @       @      �?      "@                               @                      �?      �?                              �?                      �?                                              @       @                      @                                       @      �?                      @      �?                      �?      �?                                                      �?                              @              @                     �@@      K@     @R@     @R@      @      @      @              @      @                      �?                              @      @                              @                      @      @                      @                                      @                                      @              =@     �G@      Q@     @R@      =@     �G@      P@      .@      <@     �D@     �L@      @      5@     �B@      C@       @      $@      0@      @              "@      0@      @              @      @      @              @                              @      @      @              @      @                              @                      @                                       @      @                              @                       @                       @      $@                      �?                              �?      $@                      �?       @                      �?                                       @                               @                      �?              @              �?                                              @              &@      5@      ?@       @      &@      5@      9@       @      �?      �?      $@                      �?      $@                      �?      @                              @                      �?       @                      �?                                       @                              @              �?                              $@      4@      .@       @      @      &@      �?              �?      &@      �?              �?      &@                              &@                      �?                                              �?              @                              @      "@      ,@       @              "@      ,@       @              "@      �?                              �?                      "@                                      *@       @                      (@                              �?       @                              �?                      �?      �?                      �?                                      �?      @                                              @              @      @      3@       @      @              .@               @                              @              .@               @                               @              .@                              "@               @              @               @                                              @              �?      @      @       @               @               @               @                                               @      �?       @      @              �?       @                              �?                      �?      �?                      �?                                      �?                                      @              �?      @      @      &@               @      �?      $@               @      �?                       @                                      �?                                      $@      �?      @      @      �?              @              �?              @                                              �?      �?              @              �?                                              @                              @      M@                      @      9@                              ,@                      @      &@                              &@                      @                                     �@@      A@      0@      3@      ,@      @@      @                              @                      @@                               @      *@      3@      ,@       @       @      @      @       @      �?      @      �?                              �?       @      �?      @               @      �?      �?                              �?               @      �?                       @                                      �?                                      @                      @              @               @              @               @              �?               @                                              �?                               @              @                              @      .@      $@              @      �?       @              @                                      �?       @                      �?      �?                              �?                      �?                                      �?              �?      ,@       @                      "@                      �?      @       @              �?      @                              @                      �?      �?                              �?                      �?                                               @      �?              �?       @      �?                                              �?       @                      �?                                       @�t�bub�V�      hhubh)��}�(hhhhhNhKhKhG        hh$hNhJg}�XhG        hNhG        hHKhIKhJh(h+K ��h-��R�(KK��hb�C               �?       @      @�t�bhVhghQC       ���R�hkKhlhoKh(h+K ��h-��R�(KK��hQ�C       �t�bK��R�}�(hKhyM�hzh(h+K ��h-��R�(KM���h��B��         �                   �@������?�            �@       �                    �?��`���?           (�@              	            �@z���?1�?           @z@                          �N@hl��f�?^            �a@                           x�@�ת2�%�?]            `a@              	            ~�@�q�q�?A             X@������������������������       �        2            @Q@       	                    �? 7���B�?             ;@������������������������       �                     *@
                           @@4և���?	             ,@������������������������       �                     �?������������������������       �                     *@                           �@X�EQ]N�?            �E@������������������������       �                     �?                           �?�����?             E@������������������������       �                     2@              	            ��@r�q��?             8@                           ��@�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?                           @���Q��?             @������������������������       �                      @                           �?�q�q�?             @                           �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @       �                   �2@^��'��?�            pq@       y                    @4	 � �?�            �o@       f       	            �@������?o            �e@        W                    ��@      �?Q             ^@!       8                 ����?p�� 1a�?9            @U@"       )                   �1@&G$n��?            �B@#       $                    @�$I�$I�?             @������������������������       �                      @%       (                    �?{�G�z�?             @&       '                    !@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @*       +                    9@j�Y�H��?             >@������������������������       �                      @,       -                    �@��#��Z�?             6@������������������������       �                     @.       /                    �?�ӭ�a��?
             2@������������������������       �                     �?0       5       
             %@8߄*�u�?	             1@1       2                    @�8��8��?             (@������������������������       �                     @3       4                    @r�q��?             @������������������������       �                     �?������������������������       �                     @6       7       
             (@z�G�z�?             @������������������������       �                     �?������������������������       �                     @9       P                   �D@     @�?"             H@:       E       	            ��@أp=
��?             D@;       B                    �?.y0��k�?             :@<       =                    �?�����?             5@������������������������       �                     (@>       A                    �?�<ݚ�?             "@?       @                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @C       D                    @���Q��?             @������������������������       �                      @������������������������       �                     @F       I                    @X�Cc�?             ,@G       H                    �?      �?             @������������������������       �                     @������������������������       �                     �?J       K       
             @z�G�z�?             $@������������������������       �                      @L       M                   �>@      �?              @������������������������       �                     @N       O                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @Q       V                    @      �?              @R       S                    �?؇���X�?             @������������������������       �                     @T       U       	            x�@      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?X       _       	            ��@
��ZI�?            �A@Y       ^                 `ff�? ��WV�?             :@Z       ]                    �?�����H�?             "@[       \                    ��@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     1@`       a                    :�@�����H�?             "@������������������������       �                     @b       e                    �?      �?             @c       d       
             @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?g       x                    $@�<ݚ�?             K@h       o                    �?�z�G��?             D@i       n                    ��@8�Z$���?             *@j       m                    �?�q�q�?             @k       l       	            ��@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                     $@p       s                    ��@��}*_��?             ;@q       r                    ��@���!pc�?             &@������������������������       �                     @������������������������       �                      @t       w                    �?      �?	             0@u       v                    �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     *@������������������������       �        	             ,@z       �                   �1@x�[#���?2            �S@{       �                 ����?�9[����?/            @R@|              
            �2@�g���e�?             &@}       ~       	            j�@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @�       �                    D�@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                   @N@���D�?'             O@�       �                    0�@R3���{�?&            �N@�       �                    @�HPS!��?"             J@�       �       	            ��@     ��?             @@������������������������       �                      @�       �                    �?(;L]n�?             >@������������������������       �        
             0@�       �                    4@@4և���?             ,@�       �       
             @      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     $@�       �                    @�G�z��?             4@�       �                    �?}��7�?             &@�       �                 `ff�?      �?             @������������������������       �                     �?�       �                    @z�G�z�?             @������������������������       �                     �?������������������������       �                     @�       �                    -@�Q����?             @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                     @������������������������       �                     �?�       �       	            ��@B{	�%��?             "@������������������������       �                     �?�       �                    +@      �?              @������������������������       �                     @�       �       
             @�q�q�?             @������������������������       �                     �?�       �                    /@      �?              @������������������������       �                     �?������������������������       �                     �?�       �                    @X�<ݚ�?             "@������������������������       �                     @�       �                 @33�?�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?�       �                    H@�q�q�?             @������������������������       �                     @������������������������       �                      @�       �       
             $@R�}e�.�?             :@�       �                    �?@4և���?             ,@�       �                    @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     &@�       �                    @      �?             (@������������������������       �                     @�       �                   �J@      �?              @�       �                    �?؇���X�?             @�       �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                     �?�       /                   �?��+����?           z@�       �                    �@�>�r�?y            �h@�       �                    �?g\�5�?             :@�       �       	            9�@�X�C�?             ,@�       �       
             *@����X�?             @������������������������       �                     @������������������������       �                      @������������������������       �                     @�       �       	            G�@�q�q�?	             (@������������������������       �                      @������������������������       �                     @�                          ��@:*G���?i            �e@�                          ��@&�*�¥�?W             a@�       �                   �0@�k�Vt��?J            @]@�       �                    @��a�2�?9            �T@�       �                    l�@$I�$I��?             E@�       �                    $@�m۶m��?             ,@�       �                     @�C��2(�?             &@������������������������       �                     �?������������������������       �                     $@�       �                 033�?�q�q�?             @������������������������       �                      @������������������������       �                     �?�       �       	            5�@:/����?             <@�       �       	            r�@��S���?             .@������������������������       �                      @������������������������       �                     @�       �                 ����?$�q-�?             *@������������������������       �                     @�       �                    J@؇���X�?             @������������������������       �                     �?������������������������       �                     @�       �                    �?z3�Vf`�?            �D@������������������������       �                     @�       �                 ����?�3�R��?             C@�       �                    *@$I�$I��?             ,@�       �       
            �0@�q�q�?	             (@�       �                    ��@B{	�%��?             "@������������������������       �                     �?�       �                    ,�@      �?              @������������������������       �                     @�       �                    !@      �?             @������������������������       �                     @������������������������       �                     �?�       �                    �?VUUUUU�?             @������������������������       �                     �?�       �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�       �                    @��8��8�?             8@�       �       	            @�@6�80\��?             3@������������������������       �                     @�       �                    )@�Q����?             .@�       �       
            �1@��!pc�?	             &@�       �       	            p�@ףp=
�?             $@������������������������       �                     @�       �                    4@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�       �                    �?      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�             	            �@|�l�]�?             A@�             
             3@;n,�R�?             6@�                          �?f�t���?
             1@             	            9�@���k���?             &@                        �1@�<ݚ�?             "@������������������������       �                     �?                         @      �?              @                         3@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     @������������������������       �                      @	      
                hff�?r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @                        �C@�8��8��?             (@            
             )@z�G�z�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                     @                         7@>
ףp=�?             4@������������������������       �                     @                         @�@6�h$��?	             .@������������������������       �                     &@                         T�@      �?             @������������������������       �                     �?                         @�q�q�?             @������������������������       �                      @������������������������       �                     �?                         @ȫz���?            �A@������������������������       �                     @      *                   ��@     p�?             @@      %                   �?ˠT�x�?             6@      "                  �6@�n���?             "@       !      
             )@�q�q�?             @������������������������       �                      @������������������������       �                     �?#      $                   n�@�q�q�?             @������������������������       �                     @������������������������       �                      @&      '                   �?.y0��k�?	             *@������������������������       �                     �?(      )                033@�8��8��?             (@������������������������       �                     &@������������������������       �                     �?+      ,                   @      �?             $@������������������������       �                     @-      .                   C@r�q��?             @������������������������       �                     @������������������������       �                     �?0      �                033@Y����?�            `k@1      �                   @�Q�YY��?r            `g@2      K                   @���~�?d            �d@3      D                   #@�4_�g��?             F@4      C                  �E@䃞ͪ��?             9@5      B                   A@����>4�?             5@6      A      	            ��@��>4և�?             ,@7      @                   X�@      �?              @8      ?                   @�8��8��?             @9      :                ����?      �?             @������������������������       �                     �?;      <                   �?�q�q�?             @������������������������       �                     �?=      >                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                      @������������������������       �                     @������������������������       �                     @������������������������       �                     @E      J      	            ܡ@V�Lt�<�?             3@F      I                   -@��S�ۿ?             .@G      H                   T�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@������������������������       �                     @L      U                   !@�!g��?G            �^@M      N      
             !@������?             ,@������������������������       �                     @O      P      	            d�@��ˠ�?             &@������������������������       �                     @Q      T                `ff�?      �?             @R      S                   @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @V      o                   �?����dI�?@             [@W      `                   @H�o,x�?            �C@X      [                   �?t�E]t�?             &@Y      Z                   ,�@      �?             @������������������������       �                     @������������������������       �                     �?\      _                  �K@�$I�$I�?             @]      ^      	            ã@�q�q�?             @������������������������       �                      @������������������������       �                     @������������������������       �                     �?a      h      	            ��@s
^N���?             <@b      e                ����?������?             1@c      d      	            |�@      �?             @������������������������       �                     @������������������������       �                     �?f      g                  �2@$�q-�?             *@������������������������       �                     (@������������������������       �                     �?i      n      
             *@���|���?	             &@j      m      	            �@�<ݚ�?             "@k      l                  �=@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                      @p      �      	            �@^wt4O�?'            @Q@q      �      	            �@�E]t��?             F@r      �                   ��@�>����?             ;@s      v                   �?��Q��?             4@t      u                   �?ףp=
�?             $@������������������������       �                     �?������������������������       �                     "@w      |                  �L@���Q��?             $@x      y                   "@���Q��?             @������������������������       �                      @z      {      	            ��@�q�q�?             @������������������������       �                      @������������������������       �                     �?}      �                   (@z�G�z�?             @~                         @�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                      @�      �                   �?:/����?             @�      �                   X�@      �?             @������������������������       �                      @������������������������       �                      @�      �                @33�?�q�q�?             @������������������������       �                      @������������������������       �                     �?�      �                ����?�"�O�|�?             1@�      �                   �?��S�ۿ?             .@������������������������       �                      @�      �                   @؇���X�?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @�      �                   !@H%u��?             9@�      �                   -@���!pc�?             &@������������������������       �                     @������������������������       �                      @������������������������       �        	             ,@�      �                   @ܤ�[r�?             5@�      �                   �?������?
             .@�      �                   �?"pc�
�?             &@������������������������       �                     @�      �                   B@      �?             @������������������������       �                      @������������������������       �                      @�      �                   (�@      �?             @������������������������       �                      @������������������������       �                      @������������������������       �                     @�      �                   �?     `�?             @@�      �                   �?��(\���?             4@������������������������       �                     �?�      �                  @N@�lO���?             3@�      �                   �?�����H�?             2@�      �                   @�q�q�?             @������������������������       �                     �?������������������������       �                      @�      �      
             @��S�ۿ?	             .@�      �                   #@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     (@������������������������       �                     �?�      �                   ��@��8��8�?	             (@�      �                   @����X�?             @������������������������       �                     �?�      �                   I@r�q��?             @������������������������       �                     @������������������������       �                     �?�      �                   �?�Q����?             @������������������������       �                     �?�      �                   �?      �?             @������������������������       �                     @������������������������       �                     �?�      �                   &�@L��.N�?�           ؇@�      �      
            �3@�ڦ3K�?�           ��@�                         @y�%��G�?�           8�@�      �      	            I�@v;~�i�?�            `p@�      �                   b�@���H�?b            @b@�      �      	            �@�Ы܋��?J            �Z@������������������������       �                     =@�      �                   �?���xRv�?5            �S@�      �                  �0@2(&ޏ�?	             &@�      �                   �?VUUUUU�?             @�      �                   $@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �      	            ��@l�IS�?,            �P@�      �      
             @
^N��)�?             <@������������������������       �                     @�      �                   �?&%�ݒ��?             5@�      �                   �?�g���e�?             &@�      �                  �=@B{	�%��?             "@�      �                   �?؇���X�?             @������������������������       �                     @�      �                   L�@      �?              @������������������������       �                     �?������������������������       �                     �?�      �      
             ,@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �        	             $@�      �                   �?��Ha���?            �C@�      �                   1@.y0��k�?             *@�      �                `ff�?�8��8��?             (@������������������������       �                     �?������������������������       �                     &@������������������������       �                     �?�      �                `ff�? ��WV�?             :@������������������������       �                     2@�      �                  @I@      �?              @�      �                  �D@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @�      �                ����?�V��B�?            �C@�      �      
             @     ��?             @@������������������������       �                     "@�      �                   �?��{ ��?             7@�      �                  @A@p=
ףp�?             $@������������������������       �                     @�      �                   #@�q�q�?             @������������������������       �                     �?�      �                   $�@      �?              @������������������������       �                     �?������������������������       �                     �?�      �      
            �2@8�Z$���?             *@������������������������       �                     &@������������������������       �                      @�      �      	            ��@և���X�?             @������������������������       �                     @������������������������       �                     @�                         !@XB���?C             ]@�                          �?���.�6�?             G@�      �                `ff @��2(&�?             6@�      �      	            ��@�θ�?             *@������������������������       �                     �?�      �                   ��@r�q��?             (@�      �                    @�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                     "@������������������������       �                     "@������������������������       �                     8@                         ��@`����֜?'            �Q@                         �?�8��8��?             (@                          @      �?             @������������������������       �                     �?������������������������       �                     @������������������������       �                      @������������������������       �                     M@	                         @�1T����?           |@
            	            ��@�$I�$I�?             ,@������������������������       �                      @            	            �@�q�q�?             @������������������������       �                     @������������������������       �                      @      �      	            >�@o��Gz�?           0{@      U                033�?#b.��?�            Pr@      "                  �7@c�ˇ���?U            �a@                         .�@Ԇ�ݎ��?            �B@            	            ̕@�v�`��?             ?@            
             %@�C��2(�?	             &@                         (@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @                         l�@P���Q�?             4@            
             /@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     2@                      `ff�?r�q��?             @������������������������       �                     @       !                   @�q�q�?             @������������������������       �                      @������������������������       �                     �?#      0      
             @zc���?;            @Z@$      '                   ��@�	U��6�?             A@%      &      
             @���Q��?             @������������������������       �                     @������������������������       �                      @(      -                ����?�P?��2�?             =@)      ,                   Ȟ@ףp=
�?	             4@*      +      	            ��@�}�+r��?             3@������������������������       �                     2@������������������������       �                     �?������������������������       �                     �?.      /                  @H@X�<ݚ�?             "@������������������������       �                     @������������������������       �                     @1      6                   �?��.F�l�?(            �Q@2      3      
            �0@ףp=
�?             $@������������������������       �                      @4      5                   @      �?              @������������������������       �                     �?������������������������       �                     �?7      B                   @�n�E��?#            �N@8      A                  �G@j�V���?             6@9      :                   ��@�$I�$I�?
             ,@������������������������       �                     @;      >                   @j�V���?             &@<      =                   @�����H�?             "@������������������������       �                      @������������������������       �                     �??      @                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @C      N                   �?~C_j��?            �C@D      E                   p�@�>�>��?
             .@������������������������       �                     �?F      G                   @�$I�$I�?	             ,@������������������������       �                     @H      I                   `�@j�V���?             &@������������������������       �                     @J      K                   @      �?             @������������������������       �                     �?L      M                   #@�q�q�?             @������������������������       �                      @������������������������       �                     �?O      P      	            t�@      �?             8@������������������������       �                     $@Q      T                   �?      �?             ,@R      S      
             1@�<ݚ�?             "@������������������������       �                     @������������������������       �                      @������������������������       �                     @V      _      	            ��@	�i�|�?_            �b@W      X      	            Ć@$G$n��?            �B@������������������������       �                     8@Y      ^                  �J@�n_Y�K�?
             *@Z      ]      
             @z�G�z�?             $@[      \                   6�@�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     @������������������������       �                     @`      �                  �J@�mLu��?F            �\@a      p      	            M�@R.�D���?<            �W@b      m      
            �2@�?�P�a�?%             N@c      l                   �?x�}b~|�?#            �L@d      i      
             )@z�G�z�?             9@e      h                   @P���Q�?             4@f      g                  �C@r�q��?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     ,@j      k                  @C@z�G�z�?             @������������������������       �                     @������������������������       �                     �?������������������������       �                     @@n      o                   (@�q�q�?             @������������������������       �                      @������������������������       �                     �?q      z                   "@���Q��?            �A@r      s                   �?�ӭ�a��?             2@������������������������       �                     $@t      y                   p�@      �?              @u      x                   �?r�q��?             @v      w      	            �@      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                     @������������������������       �                      @{      �      	            ��@�"�O�|�?
             1@|      }                   �?�q�q�?             (@������������������������       �                      @~            	            ��@z�G�z�?             $@������������������������       �                      @������������������������       �                      @�      �                   @z�G�z�?             @������������������������       �                     @������������������������       �                     �?�      �                   @�$�_�?
             3@������������������������       �                     @�      �      
            �1@H�7�&��?             .@�      �                  �3@؇���X�?             ,@�      �                   @$�q-�?             *@������������������������       �                     �?������������������������       �                     (@������������������������       �                     �?������������������������       �                     �?�      �      	            ��@,�d�vK�?^            �a@�      �                   @��X��?             <@�      �                   |�@z�G�z�?             4@�      �                   #@�����H�?             2@�      �                   ��@      �?              @������������������������       �                     �?������������������������       �                     �?�      �                   .�@      �?	             0@������������������������       �                     *@�      �                   ,@�q�q�?             @������������������������       �                      @������������������������       �                     �?������������������������       �                      @�      �                   �?      �?              @������������������������       �                     @�      �                   ��@���Q��?             @������������������������       �                     �?�      �                   �?      �?             @�      �                   �?      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @�      �                   �?0�)AU��?L            �\@�      �                   ��@���7�?             F@������������������������       �                      @������������������������       �                     E@������������������������       �        /            �Q@�      �                `ff�?�6w)���?            �F@�      �                   '@��W���?             7@������������������������       �                      @�      �                   #@v�"���?             5@�      �                   ��@{�G�z�?
             4@�      �                   �?&���^B�?	             2@�      �                   @     ��?             0@������������������������       �                     @������������������������       �                     *@�      �                    @      �?              @������������������������       �                     �?������������������������       �                     �?������������������������       �                      @������������������������       �                     �?�      �                   &�@;n,�R�?             6@�      �                   @�������?             (@�      �                   D�@�n���?             "@�      �                   ��@և���X�?             @������������������������       �                     @�      �                  �M@      �?             @������������������������       �                     @������������������������       �                     �?������������������������       �                      @�      �                   �?�q�q�?             @������������������������       �                     �?������������������������       �                      @������������������������       �                     $@������������������������       �                     @�t�bh�h(h+K ��h-��R�(KM�KK��hb�B`X       w@     py@     �y@     �y@     �o@     `l@     `k@      a@     �a@     �\@      ]@      I@     �`@       @                     �`@      @                     �W@      �?                     @Q@                              :@      �?                      *@                              *@      �?                              �?                      *@                              C@      @                              �?                      C@      @                      2@                              4@      @                      2@      �?                      2@                                      �?                       @      @                               @                       @      �?                      �?      �?                      �?                                      �?                      �?                                       @                      @     �Z@      ]@      I@      @     �U@     @[@      I@      @     @P@      O@      E@      @     @P@      I@              @     �C@      E@               @      $@      9@              �?      @       @                       @                      �?       @       @              �?               @                               @              �?                                       @                      �?      @      7@                               @              �?      @      .@                      @                      �?       @      .@                      �?                      �?      �?      .@              �?              &@                              @              �?              @              �?                                              @                      �?      @                      �?                                      @               @      =@      1@               @      ;@      &@               @      6@       @               @      3@                              (@                       @      @                       @      �?                              �?                       @                                      @                              @       @                               @                      @                              @      "@                      @      �?                      @                                      �?                       @       @                               @                       @      @                              @                       @      �?                              �?                       @                               @      @                      �?      @                              @                      �?      @                      �?                                      @                      �?                      �?      :@       @              �?      9@                      �?       @                      �?       @                      �?                                       @                              @                              1@                              �?       @                              @                      �?      @                      �?       @                      �?                                       @                              �?                              (@      E@                      (@      <@                       @      &@                       @      �?                      �?      �?                      �?                                      �?                      �?                                      $@                      $@      1@                       @      @                              @                       @                               @      ,@                       @      �?                              �?                       @                                      *@                              ,@       @      6@     �G@       @       @      2@     �G@      @              @      @      �?              @       @                      @                                       @                              �?      �?                      �?                                      �?       @      &@      F@      @       @      $@      F@      @       @      @      D@      @              @      =@                       @                              �?      =@                              0@                      �?      *@                      �?      @                              @                      �?                                      $@               @       @      &@      @      �?       @      @      @              �?      �?      @              �?                                      �?      @                      �?                                      @      �?      �?      @                      �?                      �?              @                              @              �?                              �?              @      �?      �?                                              @      �?                      @                               @      �?                      �?                              �?      �?                              �?                      �?                      @      @                      @                               @      @                       @                                      @                      �?                              @               @              @                                               @              3@      @                      *@      �?                       @      �?                              �?                       @                              &@                              @      @                              @                      @       @                      @      �?                       @      �?                       @                                      �?                      @                                      �?             �\@     @\@     �Y@     �U@      Q@      K@     �E@     �@@      *@       @      &@              @       @      @              @       @                      @                                       @                                      @               @              @               @                                              @             �K@      J@      @@     �@@     �A@     �F@      9@      @@      A@      C@      8@      5@      ;@      9@      5@      $@      3@      $@      *@              &@       @      �?              $@              �?                              �?              $@                              �?       @                               @                      �?                               @       @      (@               @      @                       @                                      @                              �?      (@                              @                      �?      @                      �?                                      @               @      .@       @      $@                      @               @      .@      @      $@      @      �?       @      @       @      �?       @      @      �?              �?      @                      �?              �?                      @                              @      �?                      @                              @      �?                              �?      �?      �?              �?                                      �?      �?                      �?                                      �?               @                              @      ,@      @      @      @      "@      @      @      @                                      "@      @      @              "@      �?      �?              "@      �?                      @                               @      �?                              �?                       @                                              �?                       @       @                       @                                       @              @                      @      *@      @      &@      @      *@       @              @       @       @               @      @       @               @      @                      �?                              �?      @                      �?       @                               @                      �?                                      @                                       @              @      �?                      @                                      �?                              @                                      �?      &@                      �?      @                      �?                                      @                              @      �?      @      �?      &@              @                      �?       @      �?      &@                              &@      �?       @      �?              �?                                       @      �?                       @                                      �?              4@      @      @      �?                      @              4@      @      @      �?      .@       @      @      �?      @       @      @                       @      �?                       @                                      �?              @               @              @                                               @              &@              �?      �?                              �?      &@              �?              &@                                              �?              @      @                              @                      @      �?                      @                                      �?                      G@     �M@      N@      K@     �C@      M@     �D@     �H@      <@      K@     �A@     �H@      @      7@      @      $@      @      "@      @      $@      @      "@      @      @      @       @      @      @      @       @      @              @       @      �?              �?       @      �?                              �?              �?       @                              �?                      �?      �?                      �?                                      �?                       @                                               @                                      @              @                                              @      �?      ,@      @              �?      ,@                      �?       @                      �?                                       @                              (@                                      @              8@      ?@      <@     �C@       @      �?      @      �?      @                              @      �?      @      �?      @                                      �?      @      �?              �?              �?              �?                                              �?                      @              0@      >@      8@      C@      @      ,@      @      ,@       @      �?      �?      @              �?              @                              @              �?                       @              �?      @       @                      @       @                                                      @                      �?              @      *@      @      @      @      *@                      @      �?                      @                                      �?                      �?      (@                              (@                      �?                                              @      @                       @      @                       @      �?                              �?                       @                                      @                       @              $@      0@      3@      8@      $@      0@      0@       @      $@      .@       @              @      *@                      �?      "@                      �?                                      "@                      @      @                       @      @                               @                       @      �?                       @                                      �?                      @      �?                       @      �?                              �?                       @                               @                              @       @       @               @       @                       @                                       @                      �?               @                               @              �?                                      �?      ,@       @              �?      ,@                               @                      �?      @                      �?                                      @                                       @                      @      6@                      @       @                      @                                       @                              ,@      &@      @      @              &@      @                      "@       @                      @                               @       @                       @                                       @                       @       @                       @                                       @                                      @              @      �?      3@      @       @              0@       @                              �?       @              0@      �?       @              0@              �?               @              �?                                               @              �?              ,@              �?               @              �?                                               @                              (@                                      �?      @      �?      @      @      @               @                              �?              @              �?              @                                              �?                      �?      �?      @              �?                                      �?      @                              @                      �?             �\@     �f@     `h@     q@     �\@     �f@     �g@     q@     �[@      d@     �f@     0p@      B@      L@      L@     �\@      B@      L@      J@       @      ?@      A@      D@       @      =@                               @      A@      D@       @      �?       @      �?      �?      �?              �?      �?      �?                      �?                              �?      �?                                              �?                       @                      �?      :@     �C@      �?      �?      8@      @                      @                      �?      1@      @              �?      @      @              �?      @      �?              �?      @                              @                      �?      �?                              �?                      �?                                      �?      �?                      �?                                      �?                               @                      $@                               @      B@      �?              �?      &@      �?                      &@      �?                              �?                      &@                      �?                              �?      9@                              2@                      �?      @                      �?      �?                              �?                      �?                                      @              @      6@      (@              �?      6@      "@                      "@                      �?      *@      "@              �?       @      @                              @              �?       @                              �?                      �?      �?                      �?                                      �?                              &@       @                      &@                                       @              @              @              @                                              @                              @      \@                      @     �E@                      @      3@                      @      $@                      �?                               @      $@                       @      �?                       @                                      �?                              "@                              "@                              8@                      �?     @Q@                      �?      &@                      �?      @                      �?                                      @                               @                              M@     �R@      Z@     @_@      b@       @              @       @       @                                              @       @                      @                                       @     �P@      Z@     @^@     �a@     �P@      Z@     �[@      (@      A@     �B@     �P@      @      �?      0@      4@              �?      &@      3@              �?      $@                      �?       @                               @                      �?                                       @                              �?      3@                      �?      �?                      �?                                      �?                              2@                      @      �?                      @                               @      �?                       @                                      �?             �@@      5@     �G@      @      4@      @      @               @              @                              @               @                              2@      @      @              2@       @                      2@      �?                      2@                                      �?                              �?                              @      @                              @                      @                      *@      ,@      D@      @              �?      "@                               @                      �?      �?                              �?                      �?                      *@      *@      ?@      @       @      @      0@               @      @       @                      @                       @      �?       @              �?               @                               @              �?                              �?      �?                      �?                                      �?                                       @              &@      "@      .@      @      �?       @       @      @      �?                                       @       @      @                              @               @       @      �?                      @                       @      �?      �?                      �?                       @              �?               @                                              �?      $@      @      @              $@                                      @      @                       @      @                              @                       @                              @                     �@@     �P@     �E@       @      @@      @                      8@                               @      @                       @       @                      �?       @                      �?                                       @                      @                                      @                      �?      O@     �E@       @              M@      ?@      @             �J@      @                      J@      @                      4@      @                      3@      �?                      @      �?                      @                                      �?                      ,@                              �?      @                              @                      �?                              @@                              �?       @                               @                      �?                              @      8@      @              �?      .@       @                      $@                      �?      @       @              �?      @                      �?      �?                      �?                                      �?                              @                                       @              @      "@      @              @       @                       @                               @       @                       @                                       @                              �?      @                              @                      �?              �?      @      (@       @              @                      �?              (@       @                      (@       @                      (@      �?                              �?                      (@                                      �?      �?                                              &@     ``@                      "@      3@                      @      0@                       @      0@                      �?      �?                      �?                                      �?                      �?      .@                              *@                      �?       @                               @                      �?                               @                              @      @                      @                               @      @                      �?                              �?      @                      �?      �?                              �?                      �?                                       @                       @      \@                       @      E@                       @                                      E@                             �Q@      @      4@      @      ,@      �?      @      @      *@               @                      �?      @      @      *@              @      @      *@              @      �?      *@              @              *@              @                                              *@              �?      �?                              �?                      �?                                       @              �?                              @      ,@      @      �?      @      @      @      �?      @      @       @              @      @                              @                      @      �?                      @                                      �?                                       @                               @      �?                              �?                       @                      $@                                      @        �t�bubhhubehhub.